module vga_pic(
input wire vga_clk , 
input wire sys_rst_n , 
input wire [9:0] pix_x , 
input wire [9:0] pix_y , 

output reg [15:0] pix_data 

);


parameter CHAR_B_H= 10'd100 , 
CHAR_B_V= 10'd100 ; 

parameter CHAR_W = 10'd256 , 
CHAR_H = 10'd64 ; 

parameter BLACK = 16'h0000, 
WHITE = 16'hFFFF, 
GOLDEN = 16'hFEC0; 


wire [9:0] char_x ; 
wire [9:0] char_y ; 


reg [255:0] char [63:0] ; 


assign char_x = (((pix_x >= CHAR_B_H) && (pix_x < (CHAR_B_H + CHAR_W)))
&&((pix_y >= CHAR_B_V)&&(pix_y < (CHAR_B_V + CHAR_H))))
? (pix_x - CHAR_B_H) : 10'h3FF;
assign char_y = (((pix_x >= CHAR_B_H) && (pix_x < (CHAR_B_H + CHAR_W)))
&&((pix_y >= CHAR_B_V)&&(pix_y < (CHAR_B_V + CHAR_H))))
? (pix_y - CHAR_B_V) : 10'h3FF;


always@(posedge vga_clk)
begin
char[0] <= 256'h0000000000000000000000ffff0301010101010101010101010101010101010101010101010101010101010101010101010101010f7f7f000000000000000000;
char[1] <= 256'h0000000000000000000000ffffffffffffffffffffffefefefe7e7e3e3e1e1e0e0e0e0e0e0e0e0e0e0e0e0e0e0e0e0e0e0e0e0f0fcffff000000000000000000; 
char[2] <= 256'h00000000000000000000008080c0c0c0e0e0f0f0f8f8f8fcfcfefeffffffffffff7f7f7f3f3f1f1f0f0f07070303030101000000008080000000000000000000;
char[3] <= 256'h0000000000000000000000000000000000000000000000000000000000808080c0c0e0e0f0f0f8f8f8fdfdffffffffffffffff7f7f3e3e000000000000000000;
char[4] <= 256'h0000000000000000000000000000000000000000000000000101030307070f0f1f1f1f3f3e7e7cfcfcf8f8f0f0e0e0c0c0808000000000000000000000000000;
char[5] <= 256'h000000000000000000000007070f0f1f1f1f3f3f7f7ffdfdf9f9f1f1e1e1c1c181810101010101010101010101010101010101010fffff000000000000000000;
char[6] <= 256'h0000000000000000000000ffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffff000000000000000000;
char[7] <= 256'h0000000000000000000000fefec08080808080808080808080808080808080808080808080808080808080808080808080808080f0fefe000000000000000000;
char[8] <= 256'h00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
char[9] <= 256'h00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
char[10] <= 256'h00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
char[11] <= 256'h00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
char[12] <= 256'h00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
char[13] <= 256'h00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
char[14] <= 256'h00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
char[15] <= 256'h00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
char[16] <= 256'h00000000000000000000007f7f000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
char[17] <= 256'h0000000000000000000000ffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffff7f7f3f3f1f07010000000000000000000000;
char[18] <= 256'h0000000000000000000000ffffe0c0c0c0c0c0c0c0c0c0c0c0c0c0c0c0c0c0c0c0c0c0c0c0c0c0c0c0c0c0c0c0c0c0c0e0f0f8ffff1f00000000000000000000;
char[19] <= 256'h00000000000000000000008080000000000000000000000000000000000000000000000000000000000000000000000000000000feffff000000000000000000;
char[20] <= 256'h000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000003ffffe000000000000000000;
char[21] <= 256'h00000000000000000000003f3f000000000000000000000000000000000000000000000000000000000000000000000001030f7ffce000000000000000000000;
char[22] <= 256'h0000000000000000000000ffff7e3c3c3c3c3c3c3c3c3c3c3c3c3c3c3c3c3c3c3c3c3c3c3c3c3c3c3c3c3c3c3c7c7cf8f8f0c080000000000000000000000000;
char[23] <= 256'h0000000000000000000000fcfc000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
char[24] <= 256'h00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
char[25] <= 256'h00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
char[26] <= 256'h00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
char[27] <= 256'h00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
char[28] <= 256'h00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
char[29] <= 256'h00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
char[30] <= 256'h00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
char[31] <= 256'h00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
char[32] <= 256'h00000000000000000000000000000000000103030303030303010000000000000000000000000000000007070703030301010100000000000000000000000000;
char[33] <= 256'h000000000000000000000000030f3f7ffffefcfcfcfcfcfeffffff7f1f07000000000000000000000000c0c0e0f0f8fcfefffffffffc60000000000000000000;
char[34] <= 256'h00000000000000000000037ffff8c080000000000000000080e0feffffffff0f000000000000000000000000000000000080f0feff0f00000000000000000000;
char[35] <= 256'h00000000000000000000fffff10000000000000000000000000000c0fcffffffff0f000000000000000000000000000000000000feff7f000000000000000000;
char[36] <= 256'h00000000000000000000fcffff01000000000000000000000000000000e0feffffffff0f000000000000000000000000000000003fffff000000000000000000;
char[37] <= 256'h0000000000000000000000f0ffff3f0f070300000000000000000000000000e0fcffffffff3f0f03010000000000000103070f7ffffc00000000000000000000;
char[38] <= 256'h000000000000000000003078f8f8f8f8fcfcfc7c7c00000000000000000000000080e0f0fcfeffffffff7f7f7ffffffffefcf0e0800000000000000000000000;
char[39] <= 256'h00000000000000000000000000000000000000000000000000000000000000000000000000000000808080808080000000000000000000000000000000000000;
char[40] <= 256'h00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
char[41] <= 256'h00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
char[42] <= 256'h00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
char[43] <= 256'h00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
char[44] <= 256'h00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
char[45] <= 256'h00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
char[46] <= 256'h00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
char[47] <= 256'h00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
char[48] <= 256'h000000000000000000000001030307070f0f1f1f1f00000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
char[49] <= 256'h0000000000000000000000fffffff8f0e0c080000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
char[50] <= 256'h0000000000000000000000ffff000000000000000000000000000000000000000000000000000000000000000000000000000000003f3f000000000000000000;
char[51] <= 256'h0000000000000000000000ffff1f1f1f1f1f1f1f1f1f1f1f1f1f1f1f1f1f1f1f1f1f1f1f1f1f1f1f1f1f1f1f1f1f1f1f1f1f1f3fffffff000000000000000000;
char[52] <= 256'h0000000000000000000000fffff0f0f0f0f0f0f0f0f0f0f0f0f0f0f0f0f0f0f0f0f0f0f0f0f0f0f0f0f0f0f0f0f0f0f0f0f0f0f8feffff000000000000000000;
char[53] <= 256'h0000000000000000000000ffff00000000000000000000000000000000000000000000000000000000000000000000000000000000f8f8000000000000000000;
char[54] <= 256'h0000000000000000000000ffffff3f0f070303010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
char[55] <= 256'h0000000000000000000000808080c0c0e0e0f0f0f000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
char[56] <= 256'h00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
char[57] <= 256'h00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
char[58] <= 256'h00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
char[59] <= 256'h00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
char[60] <= 256'h00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
char[61] <= 256'h00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
char[62] <= 256'h00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
char[63] <= 256'h00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;

 end


 always@(posedge vga_clk or negedge sys_rst_n)
 if(sys_rst_n == 1'b0)
 pix_data <= BLACK;
 else if((((pix_x >= (CHAR_B_H - 1'b1))
 && (pix_x < (CHAR_B_H + CHAR_W -1'b1)))
 && ((pix_y >= CHAR_B_V) && (pix_y < (CHAR_B_V + CHAR_H))))
 && (char[char_y][10'd255 - char_x] == 1'b1))
 pix_data <= GOLDEN;
 else
 pix_data <= BLACK;

 endmodule
