module vga_pic(
input wire vga_clk , 
input wire sys_rst_n , 
input wire [9:0] pix_x , 
input wire [9:0] pix_y , 

output reg [15:0] pix_data 

);


//parameter define
parameter CHAR_B_H= 10'd192 , 
CHAR_B_V= 10'd208 ; 

parameter CHAR_W = 10'd256 , 
CHAR_H = 10'd64 ; 

parameter BLACK = 16'h0000, 
WHITE = 16'hFFFF, 
GOLDEN = 16'hFEC0; 

//wire define
wire [9:0] char_x ; 
wire [9:0] char_y ; 

//reg define
reg [255:0] char [63:0] ; 

////
//\* Main Code \//
////


assign char_x = (((pix_x >= CHAR_B_H) && (pix_x < (CHAR_B_H + CHAR_W)))
&&((pix_y >= CHAR_B_V)&&(pix_y < (CHAR_B_V + CHAR_H))))
? (pix_x - CHAR_B_H) : 10'h3FF;
assign char_y = (((pix_x >= CHAR_B_H) && (pix_x < (CHAR_B_H + CHAR_W)))
&&((pix_y >= CHAR_B_V)&&(pix_y < (CHAR_B_V + CHAR_H))))
? (pix_y - CHAR_B_V) : 10'h3FF;

always@(posedge vga_clk)
begin
char[0] <=  256'h0000000000000000000000000000000000000000000000000000000000000000;
char[1] <=  256'h0000000000000000000000000000000000000000000000000000000000000000;
char[2] <=  256'h0000000000000000000000000000000000000000000000000000000000000000;
char[3] <=  256'h0000000000000000000000000000000000000000000000000000000000000000;
char[4] <=  256'h0000000000000000000000000000000000000000000000000000000000000000;
char[5] <=  256'h0000000000000000000000000000000000000000000000000000000000000000;
char[6] <=  256'h0000000000000000000000000000000000000000000000000000000000000000;
char[7] <=  256'h0000000000000000000000000000000000000000000000000000000000000000;
char[8] <=  256'h0000000000000000000000000000000000000000000000000000000000000000;
char[9] <=  256'hE0FF030000E0FF070000000000000000000000FC0F0000000000000000000000;
char[10] <= 256'hF0FF070000F0FF07C0FFFF0100FCFF010000F0FFFF83010000F8FFFFFFFF1F00;
char[11] <= 256'h00FF070000F8FF0000F80F0000800F0000003E00E0FF010000FC07F007E01F00;
char[12] <= 256'h00FC0F0000F83F0000F00700000007000080070000FE0300007C00F007003F00;
char[13] <= 256'h00FC0F0000FC3F0000F007000000070000E0030000F80300003E00F007003C00;
char[14] <= 256'h00FC0F0000FC3F0000F007000000070000F0010000F00300001E00F007007800;
char[15] <= 256'h00FC1F0000FE3F0000F007000000070000F8000000E00300000F00F007007000;
char[16] <= 256'h00FC1F0000FE3F0000F007000000070000FC000000800300000700F007007000;
char[17] <= 256'h00FC3F0000FF3F0000F0070000000700007C000000000700800300F00700E000;
char[18] <= 256'h00FC3F0000EF3F0000F0070000000700007C000000000300000000F007000000;
char[19] <= 256'h00BC7F0080EF3F0000F007000000070000FC000000000000000000F007000000;
char[20] <= 256'h00BC7F0080E73F0000F007000000070000FC000000000000000000F007000000;
char[21] <= 256'h003C7F00C0E73F0000F007000000070000FC030000000000000000F007000000;
char[22] <= 256'h003CFF00C0E73F0000F007000000070000F80F0000000000000000F007000000;
char[23] <= 256'h003CFE00C0E33F0000F007000000070000F07F0000000000000000F007000000;
char[24] <= 256'h003CFE01E0E33F0000F007000000070000C0FF0700000000000000F007000000;
char[25] <= 256'h003CFE01E0E13F0000F00700000007000000FF7F00000000000000F007000000;
char[26] <= 256'h003CFC03F0E13F0000F00700000007000000F0FF07000000000000F007000000;
char[27] <= 256'h003CFC03F0E03F0000F0070000000700000080FFFF000000000000F007000000;
char[28] <= 256'h003CF803F8E03F0000F0070000000700000000F8FF070000000000F007000000;
char[29] <= 256'h003CF80778E03F0000F007000000070000000000FF3F0000000000F007000000;
char[30] <= 256'h003CF0077CE03F0000F007000000070000000000F0FF0000000000F007000000;
char[31] <= 256'h003CF00F3CE03F0000F00700000007000000000080FF0300000000F007000000;
char[32] <= 256'h003CF00F3EE03F0000F00700000007000000000000FC0700000000F007000000;
char[33] <= 256'h003CE01F1EE03F0000F00700000007000000000000F00F00000000F007000000;
char[34] <= 256'h003CE01F1FE03F0000F00700000007000000000000E01F00000000F007000000;
char[35] <= 256'h003CC01F0FE03F0000F00700000007000000000000C01F00000000F007000000;
char[36] <= 256'h003CC03F0FE03F0000F00700000007000000000000801F00000000F007000000;
char[37] <= 256'h003C80BF0FE03F0000F0070000000700000E000000801F00000000F007000000;
char[38] <= 256'h003C80FF07E03F0000F0070000000700001E000000801F00000000F007000000;
char[39] <= 256'h003C00FF07E03F0000F0070000000700003C000000801F00000000F007000000;
char[40] <= 256'h003C00FF03E03F0000F0070000000300007C000000801F00000000F007000000;
char[41] <= 256'h003C00FF03E03F0000E00F000080030000FC000000C00F00000000F007000000;
char[42] <= 256'h003C00FE01E03F0000E00F0000C0010000F8010000E00700000000F007000000;
char[43] <= 256'h003C00FE01E03F0000C01F0000F0000000F8070000F00300000000F007000000;
char[44] <= 256'h003C00FC00E03F0000007F00003E000000F83F0000FC0000000000F007000000;
char[45] <= 256'hE0FF07FC00FFFF070000FC07E00F000000F0FF03803F0000000000F81F000000;
char[46] <= 256'hE0FF077880FFFF070000C0FFFF010000007080FFFF0700000000F0FFFF070000;
char[47] <= 256'hE0FF073000FFFF07000000E003000000000000C0070000000000000000000000;
char[48] <= 256'h0000000000000000000000000000000000000000000000000000000000000000;
char[49] <= 256'h0000000000000000000000000000000000000000000000000000000000000000;
char[50] <= 256'h0000000000000000000000000000000000000000000000000000000000000000;
char[51] <= 256'h0000000000000000000000000000000000000000000000000000000000000000;
char[52] <= 256'h0000000000000000000000000000000000000000000000000000000000000000;
char[53] <= 256'h0000000000000000000000000000000000000000000000000000000000000000;
char[54] <= 256'h0000000000000000000000000000000000000000000000000000000000000000;
char[55] <= 256'h0000000000000000000000000000000000000000000000000000000000000000;
char[56] <= 256'h0000000000000000000000000000000000000000000000000000000000000000;
char[57] <= 256'h0000000000000000000000000000000000000000000000000000000000000000;
char[58] <= 256'h0000000000000000000000000000000000000000000000000000000000000000;
char[59] <= 256'h0000000000000000000000000000000000000000000000000000000000000000;
char[60] <= 256'h0000000000000000000000000000000000000000000000000000000000000000;
char[61] <= 256'h0000000000000000000000000000000000000000000000000000000000000000;
char[62] <= 256'h0000000000000000000000000000000000000000000000000000000000000000;
char[63] <= 256'h0000000000000000000000000000000000000000000000000000000000000000;
 end

 always@(posedge vga_clk or negedge sys_rst_n)
 if(sys_rst_n == 1'b0)
 pix_data <= BLACK;
 else if((((pix_x >= (CHAR_B_H - 1'b1))
 && (pix_x < (CHAR_B_H + CHAR_W -1'b1)))
 && ((pix_y >= CHAR_B_V) && (pix_y < (CHAR_B_V + CHAR_H))))
 && (char[char_y][10'd255 - char_x] == 1'b1))
 pix_data <= GOLDEN;
 else
 pix_data <= BLACK;

 endmodule
