module rom_go (clock, address, q);
input clock;
output [0:0] q;
input [14:0] address;
reg [0:0] dout;
reg [0:0] ram [32767:0];
assign q = dout;

initial begin
  ram[0]  = 1;
  ram[1]  = 1;
  ram[2]  = 1;
  ram[3]  = 1;
  ram[4]  = 1;
  ram[5]  = 1;
  ram[6]  = 1;
  ram[7]  = 1;
  ram[8]  = 1;
  ram[9]  = 1;
  ram[10]  = 1;
  ram[11]  = 1;
  ram[12]  = 1;
  ram[13]  = 1;
  ram[14]  = 1;
  ram[15]  = 1;
  ram[16]  = 1;
  ram[17]  = 1;
  ram[18]  = 1;
  ram[19]  = 1;
  ram[20]  = 1;
  ram[21]  = 1;
  ram[22]  = 1;
  ram[23]  = 1;
  ram[24]  = 1;
  ram[25]  = 1;
  ram[26]  = 1;
  ram[27]  = 1;
  ram[28]  = 1;
  ram[29]  = 1;
  ram[30]  = 1;
  ram[31]  = 1;
  ram[32]  = 1;
  ram[33]  = 1;
  ram[34]  = 1;
  ram[35]  = 1;
  ram[36]  = 1;
  ram[37]  = 1;
  ram[38]  = 1;
  ram[39]  = 1;
  ram[40]  = 1;
  ram[41]  = 1;
  ram[42]  = 1;
  ram[43]  = 1;
  ram[44]  = 1;
  ram[45]  = 1;
  ram[46]  = 1;
  ram[47]  = 1;
  ram[48]  = 1;
  ram[49]  = 1;
  ram[50]  = 1;
  ram[51]  = 1;
  ram[52]  = 1;
  ram[53]  = 1;
  ram[54]  = 1;
  ram[55]  = 1;
  ram[56]  = 1;
  ram[57]  = 1;
  ram[58]  = 1;
  ram[59]  = 1;
  ram[60]  = 1;
  ram[61]  = 1;
  ram[62]  = 1;
  ram[63]  = 1;
  ram[64]  = 1;
  ram[65]  = 1;
  ram[66]  = 1;
  ram[67]  = 1;
  ram[68]  = 1;
  ram[69]  = 1;
  ram[70]  = 1;
  ram[71]  = 1;
  ram[72]  = 1;
  ram[73]  = 1;
  ram[74]  = 1;
  ram[75]  = 1;
  ram[76]  = 1;
  ram[77]  = 1;
  ram[78]  = 1;
  ram[79]  = 1;
  ram[80]  = 1;
  ram[81]  = 1;
  ram[82]  = 1;
  ram[83]  = 1;
  ram[84]  = 1;
  ram[85]  = 1;
  ram[86]  = 1;
  ram[87]  = 1;
  ram[88]  = 1;
  ram[89]  = 1;
  ram[90]  = 1;
  ram[91]  = 1;
  ram[92]  = 1;
  ram[93]  = 1;
  ram[94]  = 1;
  ram[95]  = 1;
  ram[96]  = 1;
  ram[97]  = 1;
  ram[98]  = 1;
  ram[99]  = 1;
  ram[100]  = 1;
  ram[101]  = 1;
  ram[102]  = 1;
  ram[103]  = 1;
  ram[104]  = 1;
  ram[105]  = 1;
  ram[106]  = 1;
  ram[107]  = 1;
  ram[108]  = 1;
  ram[109]  = 1;
  ram[110]  = 1;
  ram[111]  = 1;
  ram[112]  = 1;
  ram[113]  = 1;
  ram[114]  = 1;
  ram[115]  = 1;
  ram[116]  = 1;
  ram[117]  = 1;
  ram[118]  = 1;
  ram[119]  = 1;
  ram[120]  = 1;
  ram[121]  = 1;
  ram[122]  = 1;
  ram[123]  = 1;
  ram[124]  = 1;
  ram[125]  = 1;
  ram[126]  = 1;
  ram[127]  = 1;
  ram[128]  = 1;
  ram[129]  = 1;
  ram[130]  = 1;
  ram[131]  = 1;
  ram[132]  = 1;
  ram[133]  = 1;
  ram[134]  = 1;
  ram[135]  = 1;
  ram[136]  = 1;
  ram[137]  = 1;
  ram[138]  = 1;
  ram[139]  = 1;
  ram[140]  = 1;
  ram[141]  = 1;
  ram[142]  = 1;
  ram[143]  = 1;
  ram[144]  = 1;
  ram[145]  = 1;
  ram[146]  = 1;
  ram[147]  = 1;
  ram[148]  = 1;
  ram[149]  = 1;
  ram[150]  = 1;
  ram[151]  = 1;
  ram[152]  = 1;
  ram[153]  = 1;
  ram[154]  = 1;
  ram[155]  = 1;
  ram[156]  = 1;
  ram[157]  = 1;
  ram[158]  = 1;
  ram[159]  = 1;
  ram[160]  = 1;
  ram[161]  = 1;
  ram[162]  = 1;
  ram[163]  = 1;
  ram[164]  = 1;
  ram[165]  = 1;
  ram[166]  = 1;
  ram[167]  = 1;
  ram[168]  = 1;
  ram[169]  = 1;
  ram[170]  = 1;
  ram[171]  = 1;
  ram[172]  = 1;
  ram[173]  = 1;
  ram[174]  = 1;
  ram[175]  = 1;
  ram[176]  = 1;
  ram[177]  = 1;
  ram[178]  = 1;
  ram[179]  = 1;
  ram[180]  = 1;
  ram[181]  = 1;
  ram[182]  = 1;
  ram[183]  = 1;
  ram[184]  = 1;
  ram[185]  = 1;
  ram[186]  = 1;
  ram[187]  = 1;
  ram[188]  = 1;
  ram[189]  = 1;
  ram[190]  = 1;
  ram[191]  = 1;
  ram[192]  = 1;
  ram[193]  = 1;
  ram[194]  = 1;
  ram[195]  = 1;
  ram[196]  = 1;
  ram[197]  = 1;
  ram[198]  = 1;
  ram[199]  = 1;
  ram[200]  = 1;
  ram[201]  = 1;
  ram[202]  = 1;
  ram[203]  = 1;
  ram[204]  = 1;
  ram[205]  = 1;
  ram[206]  = 1;
  ram[207]  = 1;
  ram[208]  = 1;
  ram[209]  = 1;
  ram[210]  = 1;
  ram[211]  = 1;
  ram[212]  = 1;
  ram[213]  = 1;
  ram[214]  = 1;
  ram[215]  = 1;
  ram[216]  = 1;
  ram[217]  = 1;
  ram[218]  = 1;
  ram[219]  = 1;
  ram[220]  = 1;
  ram[221]  = 1;
  ram[222]  = 1;
  ram[223]  = 1;
  ram[224]  = 1;
  ram[225]  = 1;
  ram[226]  = 1;
  ram[227]  = 1;
  ram[228]  = 1;
  ram[229]  = 1;
  ram[230]  = 1;
  ram[231]  = 1;
  ram[232]  = 1;
  ram[233]  = 1;
  ram[234]  = 1;
  ram[235]  = 1;
  ram[236]  = 1;
  ram[237]  = 1;
  ram[238]  = 1;
  ram[239]  = 1;
  ram[240]  = 1;
  ram[241]  = 1;
  ram[242]  = 1;
  ram[243]  = 1;
  ram[244]  = 1;
  ram[245]  = 1;
  ram[246]  = 1;
  ram[247]  = 1;
  ram[248]  = 1;
  ram[249]  = 1;
  ram[250]  = 1;
  ram[251]  = 1;
  ram[252]  = 1;
  ram[253]  = 1;
  ram[254]  = 1;
  ram[255]  = 1;
  ram[256]  = 1;
  ram[257]  = 1;
  ram[258]  = 1;
  ram[259]  = 1;
  ram[260]  = 1;
  ram[261]  = 1;
  ram[262]  = 1;
  ram[263]  = 1;
  ram[264]  = 1;
  ram[265]  = 1;
  ram[266]  = 1;
  ram[267]  = 1;
  ram[268]  = 1;
  ram[269]  = 1;
  ram[270]  = 1;
  ram[271]  = 1;
  ram[272]  = 1;
  ram[273]  = 1;
  ram[274]  = 1;
  ram[275]  = 1;
  ram[276]  = 1;
  ram[277]  = 1;
  ram[278]  = 1;
  ram[279]  = 1;
  ram[280]  = 1;
  ram[281]  = 1;
  ram[282]  = 1;
  ram[283]  = 1;
  ram[284]  = 1;
  ram[285]  = 1;
  ram[286]  = 1;
  ram[287]  = 1;
  ram[288]  = 1;
  ram[289]  = 1;
  ram[290]  = 1;
  ram[291]  = 1;
  ram[292]  = 1;
  ram[293]  = 1;
  ram[294]  = 1;
  ram[295]  = 1;
  ram[296]  = 1;
  ram[297]  = 1;
  ram[298]  = 1;
  ram[299]  = 1;
  ram[300]  = 1;
  ram[301]  = 1;
  ram[302]  = 1;
  ram[303]  = 1;
  ram[304]  = 1;
  ram[305]  = 1;
  ram[306]  = 1;
  ram[307]  = 1;
  ram[308]  = 1;
  ram[309]  = 1;
  ram[310]  = 1;
  ram[311]  = 1;
  ram[312]  = 1;
  ram[313]  = 1;
  ram[314]  = 1;
  ram[315]  = 1;
  ram[316]  = 1;
  ram[317]  = 1;
  ram[318]  = 1;
  ram[319]  = 1;
  ram[320]  = 1;
  ram[321]  = 1;
  ram[322]  = 1;
  ram[323]  = 1;
  ram[324]  = 1;
  ram[325]  = 1;
  ram[326]  = 1;
  ram[327]  = 1;
  ram[328]  = 1;
  ram[329]  = 1;
  ram[330]  = 1;
  ram[331]  = 1;
  ram[332]  = 1;
  ram[333]  = 1;
  ram[334]  = 1;
  ram[335]  = 1;
  ram[336]  = 1;
  ram[337]  = 1;
  ram[338]  = 1;
  ram[339]  = 1;
  ram[340]  = 1;
  ram[341]  = 1;
  ram[342]  = 1;
  ram[343]  = 1;
  ram[344]  = 1;
  ram[345]  = 1;
  ram[346]  = 1;
  ram[347]  = 1;
  ram[348]  = 1;
  ram[349]  = 1;
  ram[350]  = 1;
  ram[351]  = 1;
  ram[352]  = 1;
  ram[353]  = 1;
  ram[354]  = 1;
  ram[355]  = 1;
  ram[356]  = 1;
  ram[357]  = 1;
  ram[358]  = 1;
  ram[359]  = 1;
  ram[360]  = 1;
  ram[361]  = 1;
  ram[362]  = 1;
  ram[363]  = 1;
  ram[364]  = 1;
  ram[365]  = 1;
  ram[366]  = 1;
  ram[367]  = 1;
  ram[368]  = 1;
  ram[369]  = 1;
  ram[370]  = 1;
  ram[371]  = 1;
  ram[372]  = 1;
  ram[373]  = 1;
  ram[374]  = 1;
  ram[375]  = 1;
  ram[376]  = 1;
  ram[377]  = 1;
  ram[378]  = 1;
  ram[379]  = 1;
  ram[380]  = 1;
  ram[381]  = 1;
  ram[382]  = 1;
  ram[383]  = 1;
  ram[384]  = 1;
  ram[385]  = 1;
  ram[386]  = 1;
  ram[387]  = 1;
  ram[388]  = 1;
  ram[389]  = 1;
  ram[390]  = 1;
  ram[391]  = 1;
  ram[392]  = 1;
  ram[393]  = 1;
  ram[394]  = 1;
  ram[395]  = 1;
  ram[396]  = 1;
  ram[397]  = 1;
  ram[398]  = 1;
  ram[399]  = 1;
  ram[400]  = 1;
  ram[401]  = 1;
  ram[402]  = 1;
  ram[403]  = 1;
  ram[404]  = 1;
  ram[405]  = 1;
  ram[406]  = 1;
  ram[407]  = 1;
  ram[408]  = 1;
  ram[409]  = 1;
  ram[410]  = 1;
  ram[411]  = 1;
  ram[412]  = 1;
  ram[413]  = 1;
  ram[414]  = 1;
  ram[415]  = 1;
  ram[416]  = 1;
  ram[417]  = 1;
  ram[418]  = 1;
  ram[419]  = 1;
  ram[420]  = 1;
  ram[421]  = 1;
  ram[422]  = 1;
  ram[423]  = 1;
  ram[424]  = 1;
  ram[425]  = 1;
  ram[426]  = 1;
  ram[427]  = 1;
  ram[428]  = 1;
  ram[429]  = 1;
  ram[430]  = 1;
  ram[431]  = 1;
  ram[432]  = 1;
  ram[433]  = 1;
  ram[434]  = 1;
  ram[435]  = 1;
  ram[436]  = 1;
  ram[437]  = 1;
  ram[438]  = 1;
  ram[439]  = 1;
  ram[440]  = 1;
  ram[441]  = 1;
  ram[442]  = 1;
  ram[443]  = 1;
  ram[444]  = 1;
  ram[445]  = 1;
  ram[446]  = 1;
  ram[447]  = 1;
  ram[448]  = 1;
  ram[449]  = 1;
  ram[450]  = 1;
  ram[451]  = 1;
  ram[452]  = 1;
  ram[453]  = 1;
  ram[454]  = 1;
  ram[455]  = 1;
  ram[456]  = 1;
  ram[457]  = 1;
  ram[458]  = 1;
  ram[459]  = 1;
  ram[460]  = 1;
  ram[461]  = 1;
  ram[462]  = 1;
  ram[463]  = 1;
  ram[464]  = 1;
  ram[465]  = 1;
  ram[466]  = 1;
  ram[467]  = 1;
  ram[468]  = 1;
  ram[469]  = 1;
  ram[470]  = 1;
  ram[471]  = 1;
  ram[472]  = 1;
  ram[473]  = 1;
  ram[474]  = 1;
  ram[475]  = 1;
  ram[476]  = 1;
  ram[477]  = 1;
  ram[478]  = 1;
  ram[479]  = 1;
  ram[480]  = 1;
  ram[481]  = 1;
  ram[482]  = 1;
  ram[483]  = 1;
  ram[484]  = 1;
  ram[485]  = 1;
  ram[486]  = 1;
  ram[487]  = 1;
  ram[488]  = 1;
  ram[489]  = 1;
  ram[490]  = 1;
  ram[491]  = 1;
  ram[492]  = 1;
  ram[493]  = 1;
  ram[494]  = 1;
  ram[495]  = 1;
  ram[496]  = 1;
  ram[497]  = 1;
  ram[498]  = 1;
  ram[499]  = 1;
  ram[500]  = 1;
  ram[501]  = 1;
  ram[502]  = 1;
  ram[503]  = 1;
  ram[504]  = 1;
  ram[505]  = 1;
  ram[506]  = 1;
  ram[507]  = 1;
  ram[508]  = 1;
  ram[509]  = 1;
  ram[510]  = 1;
  ram[511]  = 1;
  ram[512]  = 1;
  ram[513]  = 1;
  ram[514]  = 1;
  ram[515]  = 1;
  ram[516]  = 1;
  ram[517]  = 1;
  ram[518]  = 1;
  ram[519]  = 1;
  ram[520]  = 1;
  ram[521]  = 1;
  ram[522]  = 1;
  ram[523]  = 1;
  ram[524]  = 1;
  ram[525]  = 1;
  ram[526]  = 1;
  ram[527]  = 1;
  ram[528]  = 1;
  ram[529]  = 1;
  ram[530]  = 1;
  ram[531]  = 1;
  ram[532]  = 1;
  ram[533]  = 1;
  ram[534]  = 1;
  ram[535]  = 1;
  ram[536]  = 1;
  ram[537]  = 1;
  ram[538]  = 1;
  ram[539]  = 1;
  ram[540]  = 1;
  ram[541]  = 1;
  ram[542]  = 1;
  ram[543]  = 1;
  ram[544]  = 1;
  ram[545]  = 1;
  ram[546]  = 1;
  ram[547]  = 1;
  ram[548]  = 1;
  ram[549]  = 1;
  ram[550]  = 1;
  ram[551]  = 1;
  ram[552]  = 1;
  ram[553]  = 1;
  ram[554]  = 1;
  ram[555]  = 1;
  ram[556]  = 1;
  ram[557]  = 1;
  ram[558]  = 1;
  ram[559]  = 1;
  ram[560]  = 1;
  ram[561]  = 1;
  ram[562]  = 1;
  ram[563]  = 1;
  ram[564]  = 1;
  ram[565]  = 1;
  ram[566]  = 1;
  ram[567]  = 1;
  ram[568]  = 1;
  ram[569]  = 1;
  ram[570]  = 1;
  ram[571]  = 1;
  ram[572]  = 1;
  ram[573]  = 1;
  ram[574]  = 1;
  ram[575]  = 1;
  ram[576]  = 1;
  ram[577]  = 1;
  ram[578]  = 1;
  ram[579]  = 1;
  ram[580]  = 1;
  ram[581]  = 1;
  ram[582]  = 1;
  ram[583]  = 1;
  ram[584]  = 1;
  ram[585]  = 1;
  ram[586]  = 1;
  ram[587]  = 1;
  ram[588]  = 1;
  ram[589]  = 1;
  ram[590]  = 1;
  ram[591]  = 1;
  ram[592]  = 1;
  ram[593]  = 1;
  ram[594]  = 1;
  ram[595]  = 1;
  ram[596]  = 1;
  ram[597]  = 1;
  ram[598]  = 1;
  ram[599]  = 1;
  ram[600]  = 1;
  ram[601]  = 1;
  ram[602]  = 1;
  ram[603]  = 1;
  ram[604]  = 1;
  ram[605]  = 1;
  ram[606]  = 1;
  ram[607]  = 1;
  ram[608]  = 1;
  ram[609]  = 1;
  ram[610]  = 1;
  ram[611]  = 1;
  ram[612]  = 1;
  ram[613]  = 1;
  ram[614]  = 1;
  ram[615]  = 1;
  ram[616]  = 1;
  ram[617]  = 1;
  ram[618]  = 1;
  ram[619]  = 1;
  ram[620]  = 1;
  ram[621]  = 1;
  ram[622]  = 1;
  ram[623]  = 1;
  ram[624]  = 1;
  ram[625]  = 1;
  ram[626]  = 1;
  ram[627]  = 1;
  ram[628]  = 1;
  ram[629]  = 1;
  ram[630]  = 1;
  ram[631]  = 1;
  ram[632]  = 1;
  ram[633]  = 1;
  ram[634]  = 1;
  ram[635]  = 1;
  ram[636]  = 1;
  ram[637]  = 1;
  ram[638]  = 1;
  ram[639]  = 1;
  ram[640]  = 1;
  ram[641]  = 1;
  ram[642]  = 1;
  ram[643]  = 1;
  ram[644]  = 1;
  ram[645]  = 1;
  ram[646]  = 1;
  ram[647]  = 1;
  ram[648]  = 1;
  ram[649]  = 1;
  ram[650]  = 1;
  ram[651]  = 1;
  ram[652]  = 1;
  ram[653]  = 1;
  ram[654]  = 1;
  ram[655]  = 1;
  ram[656]  = 1;
  ram[657]  = 1;
  ram[658]  = 1;
  ram[659]  = 1;
  ram[660]  = 1;
  ram[661]  = 1;
  ram[662]  = 1;
  ram[663]  = 1;
  ram[664]  = 1;
  ram[665]  = 1;
  ram[666]  = 1;
  ram[667]  = 1;
  ram[668]  = 1;
  ram[669]  = 1;
  ram[670]  = 1;
  ram[671]  = 1;
  ram[672]  = 1;
  ram[673]  = 1;
  ram[674]  = 1;
  ram[675]  = 1;
  ram[676]  = 1;
  ram[677]  = 1;
  ram[678]  = 1;
  ram[679]  = 1;
  ram[680]  = 1;
  ram[681]  = 1;
  ram[682]  = 1;
  ram[683]  = 1;
  ram[684]  = 1;
  ram[685]  = 1;
  ram[686]  = 1;
  ram[687]  = 1;
  ram[688]  = 1;
  ram[689]  = 1;
  ram[690]  = 1;
  ram[691]  = 1;
  ram[692]  = 1;
  ram[693]  = 1;
  ram[694]  = 1;
  ram[695]  = 1;
  ram[696]  = 1;
  ram[697]  = 1;
  ram[698]  = 1;
  ram[699]  = 1;
  ram[700]  = 1;
  ram[701]  = 1;
  ram[702]  = 1;
  ram[703]  = 1;
  ram[704]  = 1;
  ram[705]  = 1;
  ram[706]  = 1;
  ram[707]  = 1;
  ram[708]  = 1;
  ram[709]  = 1;
  ram[710]  = 1;
  ram[711]  = 1;
  ram[712]  = 1;
  ram[713]  = 1;
  ram[714]  = 1;
  ram[715]  = 1;
  ram[716]  = 1;
  ram[717]  = 1;
  ram[718]  = 1;
  ram[719]  = 1;
  ram[720]  = 1;
  ram[721]  = 1;
  ram[722]  = 1;
  ram[723]  = 1;
  ram[724]  = 1;
  ram[725]  = 1;
  ram[726]  = 1;
  ram[727]  = 1;
  ram[728]  = 1;
  ram[729]  = 1;
  ram[730]  = 1;
  ram[731]  = 1;
  ram[732]  = 1;
  ram[733]  = 1;
  ram[734]  = 1;
  ram[735]  = 1;
  ram[736]  = 1;
  ram[737]  = 1;
  ram[738]  = 1;
  ram[739]  = 1;
  ram[740]  = 1;
  ram[741]  = 1;
  ram[742]  = 1;
  ram[743]  = 1;
  ram[744]  = 1;
  ram[745]  = 1;
  ram[746]  = 1;
  ram[747]  = 1;
  ram[748]  = 1;
  ram[749]  = 1;
  ram[750]  = 1;
  ram[751]  = 1;
  ram[752]  = 1;
  ram[753]  = 1;
  ram[754]  = 1;
  ram[755]  = 1;
  ram[756]  = 1;
  ram[757]  = 1;
  ram[758]  = 1;
  ram[759]  = 1;
  ram[760]  = 1;
  ram[761]  = 1;
  ram[762]  = 1;
  ram[763]  = 1;
  ram[764]  = 1;
  ram[765]  = 1;
  ram[766]  = 1;
  ram[767]  = 1;
  ram[768]  = 1;
  ram[769]  = 1;
  ram[770]  = 1;
  ram[771]  = 1;
  ram[772]  = 1;
  ram[773]  = 1;
  ram[774]  = 1;
  ram[775]  = 1;
  ram[776]  = 1;
  ram[777]  = 1;
  ram[778]  = 1;
  ram[779]  = 1;
  ram[780]  = 1;
  ram[781]  = 1;
  ram[782]  = 1;
  ram[783]  = 1;
  ram[784]  = 1;
  ram[785]  = 1;
  ram[786]  = 1;
  ram[787]  = 1;
  ram[788]  = 1;
  ram[789]  = 1;
  ram[790]  = 1;
  ram[791]  = 1;
  ram[792]  = 1;
  ram[793]  = 1;
  ram[794]  = 1;
  ram[795]  = 1;
  ram[796]  = 1;
  ram[797]  = 1;
  ram[798]  = 1;
  ram[799]  = 1;
  ram[800]  = 1;
  ram[801]  = 1;
  ram[802]  = 1;
  ram[803]  = 1;
  ram[804]  = 1;
  ram[805]  = 1;
  ram[806]  = 1;
  ram[807]  = 1;
  ram[808]  = 1;
  ram[809]  = 1;
  ram[810]  = 1;
  ram[811]  = 1;
  ram[812]  = 1;
  ram[813]  = 1;
  ram[814]  = 1;
  ram[815]  = 1;
  ram[816]  = 1;
  ram[817]  = 1;
  ram[818]  = 1;
  ram[819]  = 1;
  ram[820]  = 1;
  ram[821]  = 1;
  ram[822]  = 1;
  ram[823]  = 1;
  ram[824]  = 1;
  ram[825]  = 1;
  ram[826]  = 1;
  ram[827]  = 1;
  ram[828]  = 1;
  ram[829]  = 1;
  ram[830]  = 1;
  ram[831]  = 1;
  ram[832]  = 1;
  ram[833]  = 1;
  ram[834]  = 1;
  ram[835]  = 1;
  ram[836]  = 1;
  ram[837]  = 1;
  ram[838]  = 1;
  ram[839]  = 1;
  ram[840]  = 1;
  ram[841]  = 1;
  ram[842]  = 1;
  ram[843]  = 1;
  ram[844]  = 1;
  ram[845]  = 1;
  ram[846]  = 1;
  ram[847]  = 1;
  ram[848]  = 1;
  ram[849]  = 1;
  ram[850]  = 1;
  ram[851]  = 1;
  ram[852]  = 1;
  ram[853]  = 1;
  ram[854]  = 1;
  ram[855]  = 1;
  ram[856]  = 1;
  ram[857]  = 1;
  ram[858]  = 1;
  ram[859]  = 1;
  ram[860]  = 1;
  ram[861]  = 1;
  ram[862]  = 1;
  ram[863]  = 1;
  ram[864]  = 1;
  ram[865]  = 1;
  ram[866]  = 1;
  ram[867]  = 1;
  ram[868]  = 1;
  ram[869]  = 1;
  ram[870]  = 1;
  ram[871]  = 1;
  ram[872]  = 1;
  ram[873]  = 1;
  ram[874]  = 1;
  ram[875]  = 1;
  ram[876]  = 1;
  ram[877]  = 1;
  ram[878]  = 1;
  ram[879]  = 1;
  ram[880]  = 1;
  ram[881]  = 1;
  ram[882]  = 1;
  ram[883]  = 1;
  ram[884]  = 1;
  ram[885]  = 1;
  ram[886]  = 1;
  ram[887]  = 1;
  ram[888]  = 1;
  ram[889]  = 1;
  ram[890]  = 1;
  ram[891]  = 1;
  ram[892]  = 1;
  ram[893]  = 1;
  ram[894]  = 1;
  ram[895]  = 1;
  ram[896]  = 1;
  ram[897]  = 1;
  ram[898]  = 1;
  ram[899]  = 1;
  ram[900]  = 1;
  ram[901]  = 1;
  ram[902]  = 1;
  ram[903]  = 1;
  ram[904]  = 1;
  ram[905]  = 1;
  ram[906]  = 1;
  ram[907]  = 1;
  ram[908]  = 1;
  ram[909]  = 1;
  ram[910]  = 1;
  ram[911]  = 1;
  ram[912]  = 1;
  ram[913]  = 1;
  ram[914]  = 1;
  ram[915]  = 1;
  ram[916]  = 1;
  ram[917]  = 1;
  ram[918]  = 1;
  ram[919]  = 1;
  ram[920]  = 1;
  ram[921]  = 1;
  ram[922]  = 1;
  ram[923]  = 1;
  ram[924]  = 1;
  ram[925]  = 1;
  ram[926]  = 1;
  ram[927]  = 1;
  ram[928]  = 1;
  ram[929]  = 1;
  ram[930]  = 1;
  ram[931]  = 1;
  ram[932]  = 1;
  ram[933]  = 1;
  ram[934]  = 1;
  ram[935]  = 1;
  ram[936]  = 1;
  ram[937]  = 1;
  ram[938]  = 1;
  ram[939]  = 1;
  ram[940]  = 1;
  ram[941]  = 1;
  ram[942]  = 1;
  ram[943]  = 1;
  ram[944]  = 1;
  ram[945]  = 1;
  ram[946]  = 1;
  ram[947]  = 1;
  ram[948]  = 1;
  ram[949]  = 1;
  ram[950]  = 1;
  ram[951]  = 1;
  ram[952]  = 1;
  ram[953]  = 1;
  ram[954]  = 1;
  ram[955]  = 1;
  ram[956]  = 1;
  ram[957]  = 1;
  ram[958]  = 1;
  ram[959]  = 1;
  ram[960]  = 1;
  ram[961]  = 1;
  ram[962]  = 1;
  ram[963]  = 1;
  ram[964]  = 1;
  ram[965]  = 1;
  ram[966]  = 1;
  ram[967]  = 1;
  ram[968]  = 1;
  ram[969]  = 1;
  ram[970]  = 1;
  ram[971]  = 1;
  ram[972]  = 1;
  ram[973]  = 1;
  ram[974]  = 1;
  ram[975]  = 1;
  ram[976]  = 1;
  ram[977]  = 1;
  ram[978]  = 1;
  ram[979]  = 1;
  ram[980]  = 1;
  ram[981]  = 1;
  ram[982]  = 1;
  ram[983]  = 1;
  ram[984]  = 1;
  ram[985]  = 1;
  ram[986]  = 1;
  ram[987]  = 1;
  ram[988]  = 1;
  ram[989]  = 1;
  ram[990]  = 1;
  ram[991]  = 1;
  ram[992]  = 1;
  ram[993]  = 1;
  ram[994]  = 1;
  ram[995]  = 1;
  ram[996]  = 1;
  ram[997]  = 1;
  ram[998]  = 1;
  ram[999]  = 1;
  ram[1000]  = 1;
  ram[1001]  = 1;
  ram[1002]  = 1;
  ram[1003]  = 1;
  ram[1004]  = 1;
  ram[1005]  = 1;
  ram[1006]  = 1;
  ram[1007]  = 1;
  ram[1008]  = 1;
  ram[1009]  = 1;
  ram[1010]  = 1;
  ram[1011]  = 1;
  ram[1012]  = 1;
  ram[1013]  = 1;
  ram[1014]  = 1;
  ram[1015]  = 1;
  ram[1016]  = 1;
  ram[1017]  = 1;
  ram[1018]  = 1;
  ram[1019]  = 1;
  ram[1020]  = 1;
  ram[1021]  = 1;
  ram[1022]  = 1;
  ram[1023]  = 1;
  ram[1024]  = 1;
  ram[1025]  = 1;
  ram[1026]  = 1;
  ram[1027]  = 1;
  ram[1028]  = 1;
  ram[1029]  = 1;
  ram[1030]  = 1;
  ram[1031]  = 1;
  ram[1032]  = 1;
  ram[1033]  = 1;
  ram[1034]  = 1;
  ram[1035]  = 1;
  ram[1036]  = 1;
  ram[1037]  = 1;
  ram[1038]  = 1;
  ram[1039]  = 1;
  ram[1040]  = 1;
  ram[1041]  = 1;
  ram[1042]  = 1;
  ram[1043]  = 1;
  ram[1044]  = 1;
  ram[1045]  = 1;
  ram[1046]  = 1;
  ram[1047]  = 1;
  ram[1048]  = 1;
  ram[1049]  = 1;
  ram[1050]  = 1;
  ram[1051]  = 1;
  ram[1052]  = 1;
  ram[1053]  = 1;
  ram[1054]  = 1;
  ram[1055]  = 1;
  ram[1056]  = 1;
  ram[1057]  = 1;
  ram[1058]  = 1;
  ram[1059]  = 1;
  ram[1060]  = 1;
  ram[1061]  = 1;
  ram[1062]  = 1;
  ram[1063]  = 1;
  ram[1064]  = 1;
  ram[1065]  = 1;
  ram[1066]  = 1;
  ram[1067]  = 1;
  ram[1068]  = 1;
  ram[1069]  = 1;
  ram[1070]  = 1;
  ram[1071]  = 1;
  ram[1072]  = 1;
  ram[1073]  = 1;
  ram[1074]  = 1;
  ram[1075]  = 1;
  ram[1076]  = 1;
  ram[1077]  = 1;
  ram[1078]  = 1;
  ram[1079]  = 1;
  ram[1080]  = 1;
  ram[1081]  = 1;
  ram[1082]  = 1;
  ram[1083]  = 1;
  ram[1084]  = 1;
  ram[1085]  = 1;
  ram[1086]  = 1;
  ram[1087]  = 1;
  ram[1088]  = 1;
  ram[1089]  = 1;
  ram[1090]  = 1;
  ram[1091]  = 1;
  ram[1092]  = 1;
  ram[1093]  = 1;
  ram[1094]  = 1;
  ram[1095]  = 1;
  ram[1096]  = 1;
  ram[1097]  = 1;
  ram[1098]  = 1;
  ram[1099]  = 1;
  ram[1100]  = 1;
  ram[1101]  = 1;
  ram[1102]  = 1;
  ram[1103]  = 1;
  ram[1104]  = 1;
  ram[1105]  = 1;
  ram[1106]  = 1;
  ram[1107]  = 1;
  ram[1108]  = 1;
  ram[1109]  = 1;
  ram[1110]  = 1;
  ram[1111]  = 1;
  ram[1112]  = 1;
  ram[1113]  = 1;
  ram[1114]  = 1;
  ram[1115]  = 1;
  ram[1116]  = 1;
  ram[1117]  = 1;
  ram[1118]  = 1;
  ram[1119]  = 1;
  ram[1120]  = 1;
  ram[1121]  = 1;
  ram[1122]  = 1;
  ram[1123]  = 1;
  ram[1124]  = 1;
  ram[1125]  = 1;
  ram[1126]  = 1;
  ram[1127]  = 1;
  ram[1128]  = 1;
  ram[1129]  = 1;
  ram[1130]  = 1;
  ram[1131]  = 1;
  ram[1132]  = 1;
  ram[1133]  = 1;
  ram[1134]  = 1;
  ram[1135]  = 1;
  ram[1136]  = 1;
  ram[1137]  = 1;
  ram[1138]  = 1;
  ram[1139]  = 1;
  ram[1140]  = 1;
  ram[1141]  = 1;
  ram[1142]  = 1;
  ram[1143]  = 1;
  ram[1144]  = 1;
  ram[1145]  = 1;
  ram[1146]  = 1;
  ram[1147]  = 1;
  ram[1148]  = 1;
  ram[1149]  = 1;
  ram[1150]  = 1;
  ram[1151]  = 1;
  ram[1152]  = 1;
  ram[1153]  = 1;
  ram[1154]  = 1;
  ram[1155]  = 1;
  ram[1156]  = 1;
  ram[1157]  = 1;
  ram[1158]  = 1;
  ram[1159]  = 1;
  ram[1160]  = 1;
  ram[1161]  = 1;
  ram[1162]  = 1;
  ram[1163]  = 1;
  ram[1164]  = 1;
  ram[1165]  = 1;
  ram[1166]  = 1;
  ram[1167]  = 1;
  ram[1168]  = 1;
  ram[1169]  = 1;
  ram[1170]  = 1;
  ram[1171]  = 1;
  ram[1172]  = 1;
  ram[1173]  = 1;
  ram[1174]  = 1;
  ram[1175]  = 1;
  ram[1176]  = 1;
  ram[1177]  = 1;
  ram[1178]  = 1;
  ram[1179]  = 1;
  ram[1180]  = 1;
  ram[1181]  = 1;
  ram[1182]  = 1;
  ram[1183]  = 1;
  ram[1184]  = 1;
  ram[1185]  = 1;
  ram[1186]  = 1;
  ram[1187]  = 1;
  ram[1188]  = 1;
  ram[1189]  = 1;
  ram[1190]  = 1;
  ram[1191]  = 1;
  ram[1192]  = 1;
  ram[1193]  = 1;
  ram[1194]  = 1;
  ram[1195]  = 1;
  ram[1196]  = 1;
  ram[1197]  = 1;
  ram[1198]  = 1;
  ram[1199]  = 1;
  ram[1200]  = 1;
  ram[1201]  = 1;
  ram[1202]  = 1;
  ram[1203]  = 1;
  ram[1204]  = 1;
  ram[1205]  = 1;
  ram[1206]  = 1;
  ram[1207]  = 1;
  ram[1208]  = 1;
  ram[1209]  = 1;
  ram[1210]  = 1;
  ram[1211]  = 1;
  ram[1212]  = 1;
  ram[1213]  = 1;
  ram[1214]  = 1;
  ram[1215]  = 1;
  ram[1216]  = 1;
  ram[1217]  = 1;
  ram[1218]  = 1;
  ram[1219]  = 1;
  ram[1220]  = 1;
  ram[1221]  = 1;
  ram[1222]  = 1;
  ram[1223]  = 1;
  ram[1224]  = 1;
  ram[1225]  = 1;
  ram[1226]  = 1;
  ram[1227]  = 1;
  ram[1228]  = 1;
  ram[1229]  = 1;
  ram[1230]  = 1;
  ram[1231]  = 1;
  ram[1232]  = 1;
  ram[1233]  = 1;
  ram[1234]  = 1;
  ram[1235]  = 1;
  ram[1236]  = 1;
  ram[1237]  = 1;
  ram[1238]  = 1;
  ram[1239]  = 1;
  ram[1240]  = 1;
  ram[1241]  = 1;
  ram[1242]  = 1;
  ram[1243]  = 1;
  ram[1244]  = 1;
  ram[1245]  = 1;
  ram[1246]  = 1;
  ram[1247]  = 1;
  ram[1248]  = 1;
  ram[1249]  = 1;
  ram[1250]  = 1;
  ram[1251]  = 1;
  ram[1252]  = 1;
  ram[1253]  = 1;
  ram[1254]  = 1;
  ram[1255]  = 1;
  ram[1256]  = 1;
  ram[1257]  = 1;
  ram[1258]  = 1;
  ram[1259]  = 1;
  ram[1260]  = 1;
  ram[1261]  = 1;
  ram[1262]  = 1;
  ram[1263]  = 1;
  ram[1264]  = 1;
  ram[1265]  = 1;
  ram[1266]  = 1;
  ram[1267]  = 1;
  ram[1268]  = 1;
  ram[1269]  = 1;
  ram[1270]  = 1;
  ram[1271]  = 1;
  ram[1272]  = 1;
  ram[1273]  = 1;
  ram[1274]  = 1;
  ram[1275]  = 1;
  ram[1276]  = 1;
  ram[1277]  = 1;
  ram[1278]  = 1;
  ram[1279]  = 1;
  ram[1280]  = 1;
  ram[1281]  = 1;
  ram[1282]  = 1;
  ram[1283]  = 1;
  ram[1284]  = 1;
  ram[1285]  = 1;
  ram[1286]  = 1;
  ram[1287]  = 1;
  ram[1288]  = 1;
  ram[1289]  = 1;
  ram[1290]  = 1;
  ram[1291]  = 1;
  ram[1292]  = 1;
  ram[1293]  = 1;
  ram[1294]  = 1;
  ram[1295]  = 1;
  ram[1296]  = 1;
  ram[1297]  = 1;
  ram[1298]  = 1;
  ram[1299]  = 1;
  ram[1300]  = 1;
  ram[1301]  = 1;
  ram[1302]  = 1;
  ram[1303]  = 1;
  ram[1304]  = 1;
  ram[1305]  = 1;
  ram[1306]  = 1;
  ram[1307]  = 1;
  ram[1308]  = 1;
  ram[1309]  = 1;
  ram[1310]  = 1;
  ram[1311]  = 1;
  ram[1312]  = 1;
  ram[1313]  = 1;
  ram[1314]  = 1;
  ram[1315]  = 1;
  ram[1316]  = 1;
  ram[1317]  = 1;
  ram[1318]  = 1;
  ram[1319]  = 1;
  ram[1320]  = 1;
  ram[1321]  = 1;
  ram[1322]  = 1;
  ram[1323]  = 1;
  ram[1324]  = 1;
  ram[1325]  = 1;
  ram[1326]  = 1;
  ram[1327]  = 1;
  ram[1328]  = 1;
  ram[1329]  = 1;
  ram[1330]  = 1;
  ram[1331]  = 1;
  ram[1332]  = 1;
  ram[1333]  = 1;
  ram[1334]  = 1;
  ram[1335]  = 1;
  ram[1336]  = 1;
  ram[1337]  = 1;
  ram[1338]  = 1;
  ram[1339]  = 1;
  ram[1340]  = 1;
  ram[1341]  = 1;
  ram[1342]  = 1;
  ram[1343]  = 1;
  ram[1344]  = 1;
  ram[1345]  = 1;
  ram[1346]  = 1;
  ram[1347]  = 1;
  ram[1348]  = 1;
  ram[1349]  = 1;
  ram[1350]  = 1;
  ram[1351]  = 1;
  ram[1352]  = 1;
  ram[1353]  = 1;
  ram[1354]  = 1;
  ram[1355]  = 1;
  ram[1356]  = 1;
  ram[1357]  = 1;
  ram[1358]  = 1;
  ram[1359]  = 1;
  ram[1360]  = 1;
  ram[1361]  = 1;
  ram[1362]  = 1;
  ram[1363]  = 1;
  ram[1364]  = 1;
  ram[1365]  = 1;
  ram[1366]  = 1;
  ram[1367]  = 1;
  ram[1368]  = 1;
  ram[1369]  = 1;
  ram[1370]  = 1;
  ram[1371]  = 1;
  ram[1372]  = 1;
  ram[1373]  = 1;
  ram[1374]  = 1;
  ram[1375]  = 1;
  ram[1376]  = 1;
  ram[1377]  = 1;
  ram[1378]  = 1;
  ram[1379]  = 1;
  ram[1380]  = 1;
  ram[1381]  = 1;
  ram[1382]  = 1;
  ram[1383]  = 1;
  ram[1384]  = 1;
  ram[1385]  = 1;
  ram[1386]  = 1;
  ram[1387]  = 1;
  ram[1388]  = 1;
  ram[1389]  = 1;
  ram[1390]  = 1;
  ram[1391]  = 1;
  ram[1392]  = 1;
  ram[1393]  = 1;
  ram[1394]  = 1;
  ram[1395]  = 1;
  ram[1396]  = 1;
  ram[1397]  = 1;
  ram[1398]  = 1;
  ram[1399]  = 1;
  ram[1400]  = 1;
  ram[1401]  = 1;
  ram[1402]  = 1;
  ram[1403]  = 1;
  ram[1404]  = 1;
  ram[1405]  = 1;
  ram[1406]  = 1;
  ram[1407]  = 1;
  ram[1408]  = 1;
  ram[1409]  = 1;
  ram[1410]  = 1;
  ram[1411]  = 1;
  ram[1412]  = 1;
  ram[1413]  = 1;
  ram[1414]  = 1;
  ram[1415]  = 1;
  ram[1416]  = 1;
  ram[1417]  = 1;
  ram[1418]  = 1;
  ram[1419]  = 1;
  ram[1420]  = 1;
  ram[1421]  = 1;
  ram[1422]  = 1;
  ram[1423]  = 1;
  ram[1424]  = 1;
  ram[1425]  = 1;
  ram[1426]  = 1;
  ram[1427]  = 1;
  ram[1428]  = 1;
  ram[1429]  = 1;
  ram[1430]  = 1;
  ram[1431]  = 1;
  ram[1432]  = 1;
  ram[1433]  = 1;
  ram[1434]  = 1;
  ram[1435]  = 1;
  ram[1436]  = 1;
  ram[1437]  = 1;
  ram[1438]  = 1;
  ram[1439]  = 1;
  ram[1440]  = 1;
  ram[1441]  = 1;
  ram[1442]  = 1;
  ram[1443]  = 1;
  ram[1444]  = 1;
  ram[1445]  = 1;
  ram[1446]  = 1;
  ram[1447]  = 1;
  ram[1448]  = 1;
  ram[1449]  = 1;
  ram[1450]  = 1;
  ram[1451]  = 1;
  ram[1452]  = 1;
  ram[1453]  = 1;
  ram[1454]  = 1;
  ram[1455]  = 1;
  ram[1456]  = 1;
  ram[1457]  = 1;
  ram[1458]  = 1;
  ram[1459]  = 1;
  ram[1460]  = 1;
  ram[1461]  = 1;
  ram[1462]  = 1;
  ram[1463]  = 1;
  ram[1464]  = 1;
  ram[1465]  = 1;
  ram[1466]  = 1;
  ram[1467]  = 1;
  ram[1468]  = 1;
  ram[1469]  = 1;
  ram[1470]  = 1;
  ram[1471]  = 1;
  ram[1472]  = 1;
  ram[1473]  = 1;
  ram[1474]  = 1;
  ram[1475]  = 1;
  ram[1476]  = 1;
  ram[1477]  = 1;
  ram[1478]  = 1;
  ram[1479]  = 1;
  ram[1480]  = 1;
  ram[1481]  = 1;
  ram[1482]  = 1;
  ram[1483]  = 1;
  ram[1484]  = 1;
  ram[1485]  = 1;
  ram[1486]  = 1;
  ram[1487]  = 1;
  ram[1488]  = 1;
  ram[1489]  = 1;
  ram[1490]  = 1;
  ram[1491]  = 1;
  ram[1492]  = 1;
  ram[1493]  = 1;
  ram[1494]  = 1;
  ram[1495]  = 1;
  ram[1496]  = 1;
  ram[1497]  = 1;
  ram[1498]  = 1;
  ram[1499]  = 1;
  ram[1500]  = 1;
  ram[1501]  = 1;
  ram[1502]  = 1;
  ram[1503]  = 1;
  ram[1504]  = 1;
  ram[1505]  = 1;
  ram[1506]  = 1;
  ram[1507]  = 1;
  ram[1508]  = 1;
  ram[1509]  = 1;
  ram[1510]  = 1;
  ram[1511]  = 1;
  ram[1512]  = 1;
  ram[1513]  = 1;
  ram[1514]  = 1;
  ram[1515]  = 1;
  ram[1516]  = 1;
  ram[1517]  = 1;
  ram[1518]  = 1;
  ram[1519]  = 1;
  ram[1520]  = 1;
  ram[1521]  = 1;
  ram[1522]  = 1;
  ram[1523]  = 1;
  ram[1524]  = 1;
  ram[1525]  = 1;
  ram[1526]  = 1;
  ram[1527]  = 1;
  ram[1528]  = 1;
  ram[1529]  = 1;
  ram[1530]  = 1;
  ram[1531]  = 1;
  ram[1532]  = 1;
  ram[1533]  = 1;
  ram[1534]  = 1;
  ram[1535]  = 1;
  ram[1536]  = 1;
  ram[1537]  = 1;
  ram[1538]  = 1;
  ram[1539]  = 1;
  ram[1540]  = 1;
  ram[1541]  = 1;
  ram[1542]  = 1;
  ram[1543]  = 1;
  ram[1544]  = 1;
  ram[1545]  = 1;
  ram[1546]  = 1;
  ram[1547]  = 1;
  ram[1548]  = 1;
  ram[1549]  = 1;
  ram[1550]  = 1;
  ram[1551]  = 1;
  ram[1552]  = 1;
  ram[1553]  = 1;
  ram[1554]  = 1;
  ram[1555]  = 1;
  ram[1556]  = 1;
  ram[1557]  = 1;
  ram[1558]  = 1;
  ram[1559]  = 1;
  ram[1560]  = 1;
  ram[1561]  = 1;
  ram[1562]  = 1;
  ram[1563]  = 1;
  ram[1564]  = 1;
  ram[1565]  = 1;
  ram[1566]  = 1;
  ram[1567]  = 1;
  ram[1568]  = 1;
  ram[1569]  = 1;
  ram[1570]  = 1;
  ram[1571]  = 1;
  ram[1572]  = 1;
  ram[1573]  = 1;
  ram[1574]  = 1;
  ram[1575]  = 1;
  ram[1576]  = 1;
  ram[1577]  = 1;
  ram[1578]  = 1;
  ram[1579]  = 1;
  ram[1580]  = 1;
  ram[1581]  = 1;
  ram[1582]  = 1;
  ram[1583]  = 1;
  ram[1584]  = 1;
  ram[1585]  = 1;
  ram[1586]  = 1;
  ram[1587]  = 1;
  ram[1588]  = 1;
  ram[1589]  = 1;
  ram[1590]  = 1;
  ram[1591]  = 1;
  ram[1592]  = 1;
  ram[1593]  = 1;
  ram[1594]  = 1;
  ram[1595]  = 1;
  ram[1596]  = 1;
  ram[1597]  = 1;
  ram[1598]  = 1;
  ram[1599]  = 1;
  ram[1600]  = 1;
  ram[1601]  = 1;
  ram[1602]  = 1;
  ram[1603]  = 1;
  ram[1604]  = 1;
  ram[1605]  = 1;
  ram[1606]  = 1;
  ram[1607]  = 1;
  ram[1608]  = 1;
  ram[1609]  = 1;
  ram[1610]  = 1;
  ram[1611]  = 1;
  ram[1612]  = 1;
  ram[1613]  = 1;
  ram[1614]  = 1;
  ram[1615]  = 1;
  ram[1616]  = 1;
  ram[1617]  = 1;
  ram[1618]  = 1;
  ram[1619]  = 1;
  ram[1620]  = 1;
  ram[1621]  = 1;
  ram[1622]  = 1;
  ram[1623]  = 1;
  ram[1624]  = 1;
  ram[1625]  = 1;
  ram[1626]  = 1;
  ram[1627]  = 1;
  ram[1628]  = 1;
  ram[1629]  = 1;
  ram[1630]  = 1;
  ram[1631]  = 1;
  ram[1632]  = 1;
  ram[1633]  = 1;
  ram[1634]  = 1;
  ram[1635]  = 1;
  ram[1636]  = 1;
  ram[1637]  = 1;
  ram[1638]  = 1;
  ram[1639]  = 1;
  ram[1640]  = 1;
  ram[1641]  = 1;
  ram[1642]  = 1;
  ram[1643]  = 1;
  ram[1644]  = 1;
  ram[1645]  = 1;
  ram[1646]  = 1;
  ram[1647]  = 1;
  ram[1648]  = 1;
  ram[1649]  = 1;
  ram[1650]  = 1;
  ram[1651]  = 1;
  ram[1652]  = 1;
  ram[1653]  = 1;
  ram[1654]  = 1;
  ram[1655]  = 1;
  ram[1656]  = 1;
  ram[1657]  = 1;
  ram[1658]  = 1;
  ram[1659]  = 1;
  ram[1660]  = 1;
  ram[1661]  = 1;
  ram[1662]  = 1;
  ram[1663]  = 1;
  ram[1664]  = 1;
  ram[1665]  = 1;
  ram[1666]  = 1;
  ram[1667]  = 1;
  ram[1668]  = 1;
  ram[1669]  = 1;
  ram[1670]  = 1;
  ram[1671]  = 1;
  ram[1672]  = 1;
  ram[1673]  = 1;
  ram[1674]  = 1;
  ram[1675]  = 1;
  ram[1676]  = 1;
  ram[1677]  = 1;
  ram[1678]  = 1;
  ram[1679]  = 1;
  ram[1680]  = 1;
  ram[1681]  = 1;
  ram[1682]  = 1;
  ram[1683]  = 1;
  ram[1684]  = 1;
  ram[1685]  = 1;
  ram[1686]  = 1;
  ram[1687]  = 1;
  ram[1688]  = 1;
  ram[1689]  = 1;
  ram[1690]  = 1;
  ram[1691]  = 1;
  ram[1692]  = 1;
  ram[1693]  = 1;
  ram[1694]  = 1;
  ram[1695]  = 1;
  ram[1696]  = 1;
  ram[1697]  = 1;
  ram[1698]  = 1;
  ram[1699]  = 1;
  ram[1700]  = 1;
  ram[1701]  = 1;
  ram[1702]  = 1;
  ram[1703]  = 1;
  ram[1704]  = 1;
  ram[1705]  = 1;
  ram[1706]  = 1;
  ram[1707]  = 1;
  ram[1708]  = 1;
  ram[1709]  = 1;
  ram[1710]  = 1;
  ram[1711]  = 1;
  ram[1712]  = 1;
  ram[1713]  = 1;
  ram[1714]  = 1;
  ram[1715]  = 1;
  ram[1716]  = 1;
  ram[1717]  = 1;
  ram[1718]  = 1;
  ram[1719]  = 1;
  ram[1720]  = 1;
  ram[1721]  = 1;
  ram[1722]  = 1;
  ram[1723]  = 1;
  ram[1724]  = 1;
  ram[1725]  = 1;
  ram[1726]  = 1;
  ram[1727]  = 1;
  ram[1728]  = 1;
  ram[1729]  = 1;
  ram[1730]  = 1;
  ram[1731]  = 1;
  ram[1732]  = 1;
  ram[1733]  = 1;
  ram[1734]  = 1;
  ram[1735]  = 1;
  ram[1736]  = 1;
  ram[1737]  = 1;
  ram[1738]  = 1;
  ram[1739]  = 1;
  ram[1740]  = 1;
  ram[1741]  = 1;
  ram[1742]  = 1;
  ram[1743]  = 1;
  ram[1744]  = 1;
  ram[1745]  = 1;
  ram[1746]  = 1;
  ram[1747]  = 1;
  ram[1748]  = 1;
  ram[1749]  = 1;
  ram[1750]  = 1;
  ram[1751]  = 1;
  ram[1752]  = 1;
  ram[1753]  = 1;
  ram[1754]  = 1;
  ram[1755]  = 1;
  ram[1756]  = 1;
  ram[1757]  = 1;
  ram[1758]  = 1;
  ram[1759]  = 1;
  ram[1760]  = 1;
  ram[1761]  = 1;
  ram[1762]  = 1;
  ram[1763]  = 1;
  ram[1764]  = 1;
  ram[1765]  = 1;
  ram[1766]  = 1;
  ram[1767]  = 1;
  ram[1768]  = 1;
  ram[1769]  = 1;
  ram[1770]  = 1;
  ram[1771]  = 1;
  ram[1772]  = 1;
  ram[1773]  = 1;
  ram[1774]  = 1;
  ram[1775]  = 1;
  ram[1776]  = 1;
  ram[1777]  = 1;
  ram[1778]  = 1;
  ram[1779]  = 1;
  ram[1780]  = 1;
  ram[1781]  = 1;
  ram[1782]  = 1;
  ram[1783]  = 1;
  ram[1784]  = 1;
  ram[1785]  = 1;
  ram[1786]  = 1;
  ram[1787]  = 1;
  ram[1788]  = 1;
  ram[1789]  = 1;
  ram[1790]  = 1;
  ram[1791]  = 1;
  ram[1792]  = 1;
  ram[1793]  = 1;
  ram[1794]  = 1;
  ram[1795]  = 1;
  ram[1796]  = 1;
  ram[1797]  = 1;
  ram[1798]  = 1;
  ram[1799]  = 1;
  ram[1800]  = 1;
  ram[1801]  = 1;
  ram[1802]  = 1;
  ram[1803]  = 1;
  ram[1804]  = 1;
  ram[1805]  = 1;
  ram[1806]  = 1;
  ram[1807]  = 1;
  ram[1808]  = 1;
  ram[1809]  = 1;
  ram[1810]  = 1;
  ram[1811]  = 1;
  ram[1812]  = 1;
  ram[1813]  = 1;
  ram[1814]  = 1;
  ram[1815]  = 1;
  ram[1816]  = 1;
  ram[1817]  = 1;
  ram[1818]  = 1;
  ram[1819]  = 1;
  ram[1820]  = 1;
  ram[1821]  = 1;
  ram[1822]  = 1;
  ram[1823]  = 1;
  ram[1824]  = 1;
  ram[1825]  = 1;
  ram[1826]  = 1;
  ram[1827]  = 1;
  ram[1828]  = 1;
  ram[1829]  = 1;
  ram[1830]  = 1;
  ram[1831]  = 1;
  ram[1832]  = 1;
  ram[1833]  = 1;
  ram[1834]  = 1;
  ram[1835]  = 1;
  ram[1836]  = 1;
  ram[1837]  = 1;
  ram[1838]  = 1;
  ram[1839]  = 1;
  ram[1840]  = 1;
  ram[1841]  = 1;
  ram[1842]  = 1;
  ram[1843]  = 1;
  ram[1844]  = 1;
  ram[1845]  = 1;
  ram[1846]  = 1;
  ram[1847]  = 1;
  ram[1848]  = 1;
  ram[1849]  = 1;
  ram[1850]  = 1;
  ram[1851]  = 1;
  ram[1852]  = 1;
  ram[1853]  = 1;
  ram[1854]  = 1;
  ram[1855]  = 1;
  ram[1856]  = 1;
  ram[1857]  = 1;
  ram[1858]  = 1;
  ram[1859]  = 1;
  ram[1860]  = 1;
  ram[1861]  = 1;
  ram[1862]  = 1;
  ram[1863]  = 1;
  ram[1864]  = 1;
  ram[1865]  = 1;
  ram[1866]  = 1;
  ram[1867]  = 1;
  ram[1868]  = 1;
  ram[1869]  = 1;
  ram[1870]  = 1;
  ram[1871]  = 1;
  ram[1872]  = 1;
  ram[1873]  = 1;
  ram[1874]  = 1;
  ram[1875]  = 1;
  ram[1876]  = 1;
  ram[1877]  = 1;
  ram[1878]  = 1;
  ram[1879]  = 1;
  ram[1880]  = 1;
  ram[1881]  = 1;
  ram[1882]  = 1;
  ram[1883]  = 1;
  ram[1884]  = 1;
  ram[1885]  = 1;
  ram[1886]  = 1;
  ram[1887]  = 1;
  ram[1888]  = 1;
  ram[1889]  = 1;
  ram[1890]  = 1;
  ram[1891]  = 1;
  ram[1892]  = 1;
  ram[1893]  = 1;
  ram[1894]  = 1;
  ram[1895]  = 1;
  ram[1896]  = 1;
  ram[1897]  = 1;
  ram[1898]  = 1;
  ram[1899]  = 1;
  ram[1900]  = 1;
  ram[1901]  = 1;
  ram[1902]  = 1;
  ram[1903]  = 1;
  ram[1904]  = 1;
  ram[1905]  = 1;
  ram[1906]  = 1;
  ram[1907]  = 1;
  ram[1908]  = 1;
  ram[1909]  = 1;
  ram[1910]  = 1;
  ram[1911]  = 1;
  ram[1912]  = 1;
  ram[1913]  = 1;
  ram[1914]  = 1;
  ram[1915]  = 1;
  ram[1916]  = 1;
  ram[1917]  = 1;
  ram[1918]  = 1;
  ram[1919]  = 1;
  ram[1920]  = 1;
  ram[1921]  = 1;
  ram[1922]  = 1;
  ram[1923]  = 1;
  ram[1924]  = 1;
  ram[1925]  = 1;
  ram[1926]  = 1;
  ram[1927]  = 1;
  ram[1928]  = 1;
  ram[1929]  = 1;
  ram[1930]  = 1;
  ram[1931]  = 1;
  ram[1932]  = 1;
  ram[1933]  = 1;
  ram[1934]  = 1;
  ram[1935]  = 1;
  ram[1936]  = 1;
  ram[1937]  = 1;
  ram[1938]  = 1;
  ram[1939]  = 1;
  ram[1940]  = 1;
  ram[1941]  = 1;
  ram[1942]  = 1;
  ram[1943]  = 1;
  ram[1944]  = 1;
  ram[1945]  = 1;
  ram[1946]  = 1;
  ram[1947]  = 1;
  ram[1948]  = 1;
  ram[1949]  = 1;
  ram[1950]  = 1;
  ram[1951]  = 1;
  ram[1952]  = 1;
  ram[1953]  = 1;
  ram[1954]  = 1;
  ram[1955]  = 1;
  ram[1956]  = 1;
  ram[1957]  = 1;
  ram[1958]  = 1;
  ram[1959]  = 1;
  ram[1960]  = 1;
  ram[1961]  = 1;
  ram[1962]  = 1;
  ram[1963]  = 1;
  ram[1964]  = 1;
  ram[1965]  = 1;
  ram[1966]  = 1;
  ram[1967]  = 1;
  ram[1968]  = 1;
  ram[1969]  = 1;
  ram[1970]  = 1;
  ram[1971]  = 1;
  ram[1972]  = 1;
  ram[1973]  = 1;
  ram[1974]  = 1;
  ram[1975]  = 1;
  ram[1976]  = 1;
  ram[1977]  = 1;
  ram[1978]  = 1;
  ram[1979]  = 1;
  ram[1980]  = 1;
  ram[1981]  = 1;
  ram[1982]  = 1;
  ram[1983]  = 1;
  ram[1984]  = 1;
  ram[1985]  = 1;
  ram[1986]  = 1;
  ram[1987]  = 1;
  ram[1988]  = 1;
  ram[1989]  = 1;
  ram[1990]  = 1;
  ram[1991]  = 1;
  ram[1992]  = 1;
  ram[1993]  = 1;
  ram[1994]  = 1;
  ram[1995]  = 1;
  ram[1996]  = 1;
  ram[1997]  = 1;
  ram[1998]  = 1;
  ram[1999]  = 1;
  ram[2000]  = 1;
  ram[2001]  = 1;
  ram[2002]  = 1;
  ram[2003]  = 1;
  ram[2004]  = 1;
  ram[2005]  = 1;
  ram[2006]  = 1;
  ram[2007]  = 1;
  ram[2008]  = 1;
  ram[2009]  = 1;
  ram[2010]  = 1;
  ram[2011]  = 1;
  ram[2012]  = 1;
  ram[2013]  = 1;
  ram[2014]  = 1;
  ram[2015]  = 1;
  ram[2016]  = 1;
  ram[2017]  = 1;
  ram[2018]  = 1;
  ram[2019]  = 1;
  ram[2020]  = 1;
  ram[2021]  = 1;
  ram[2022]  = 1;
  ram[2023]  = 1;
  ram[2024]  = 1;
  ram[2025]  = 1;
  ram[2026]  = 1;
  ram[2027]  = 1;
  ram[2028]  = 1;
  ram[2029]  = 1;
  ram[2030]  = 1;
  ram[2031]  = 1;
  ram[2032]  = 1;
  ram[2033]  = 1;
  ram[2034]  = 1;
  ram[2035]  = 1;
  ram[2036]  = 1;
  ram[2037]  = 1;
  ram[2038]  = 1;
  ram[2039]  = 1;
  ram[2040]  = 1;
  ram[2041]  = 1;
  ram[2042]  = 1;
  ram[2043]  = 1;
  ram[2044]  = 1;
  ram[2045]  = 1;
  ram[2046]  = 1;
  ram[2047]  = 1;
  ram[2048]  = 1;
  ram[2049]  = 1;
  ram[2050]  = 1;
  ram[2051]  = 1;
  ram[2052]  = 1;
  ram[2053]  = 1;
  ram[2054]  = 1;
  ram[2055]  = 1;
  ram[2056]  = 1;
  ram[2057]  = 1;
  ram[2058]  = 1;
  ram[2059]  = 1;
  ram[2060]  = 1;
  ram[2061]  = 1;
  ram[2062]  = 1;
  ram[2063]  = 1;
  ram[2064]  = 1;
  ram[2065]  = 1;
  ram[2066]  = 1;
  ram[2067]  = 1;
  ram[2068]  = 1;
  ram[2069]  = 1;
  ram[2070]  = 1;
  ram[2071]  = 1;
  ram[2072]  = 1;
  ram[2073]  = 1;
  ram[2074]  = 1;
  ram[2075]  = 1;
  ram[2076]  = 1;
  ram[2077]  = 1;
  ram[2078]  = 1;
  ram[2079]  = 1;
  ram[2080]  = 1;
  ram[2081]  = 1;
  ram[2082]  = 1;
  ram[2083]  = 1;
  ram[2084]  = 1;
  ram[2085]  = 1;
  ram[2086]  = 1;
  ram[2087]  = 1;
  ram[2088]  = 1;
  ram[2089]  = 1;
  ram[2090]  = 1;
  ram[2091]  = 1;
  ram[2092]  = 1;
  ram[2093]  = 1;
  ram[2094]  = 1;
  ram[2095]  = 1;
  ram[2096]  = 1;
  ram[2097]  = 1;
  ram[2098]  = 1;
  ram[2099]  = 1;
  ram[2100]  = 1;
  ram[2101]  = 1;
  ram[2102]  = 1;
  ram[2103]  = 1;
  ram[2104]  = 1;
  ram[2105]  = 1;
  ram[2106]  = 1;
  ram[2107]  = 1;
  ram[2108]  = 1;
  ram[2109]  = 1;
  ram[2110]  = 1;
  ram[2111]  = 1;
  ram[2112]  = 1;
  ram[2113]  = 1;
  ram[2114]  = 1;
  ram[2115]  = 1;
  ram[2116]  = 1;
  ram[2117]  = 1;
  ram[2118]  = 1;
  ram[2119]  = 1;
  ram[2120]  = 1;
  ram[2121]  = 1;
  ram[2122]  = 1;
  ram[2123]  = 1;
  ram[2124]  = 1;
  ram[2125]  = 1;
  ram[2126]  = 1;
  ram[2127]  = 1;
  ram[2128]  = 1;
  ram[2129]  = 1;
  ram[2130]  = 1;
  ram[2131]  = 1;
  ram[2132]  = 1;
  ram[2133]  = 1;
  ram[2134]  = 1;
  ram[2135]  = 1;
  ram[2136]  = 1;
  ram[2137]  = 1;
  ram[2138]  = 1;
  ram[2139]  = 1;
  ram[2140]  = 1;
  ram[2141]  = 1;
  ram[2142]  = 1;
  ram[2143]  = 1;
  ram[2144]  = 1;
  ram[2145]  = 1;
  ram[2146]  = 1;
  ram[2147]  = 1;
  ram[2148]  = 1;
  ram[2149]  = 1;
  ram[2150]  = 1;
  ram[2151]  = 1;
  ram[2152]  = 1;
  ram[2153]  = 1;
  ram[2154]  = 1;
  ram[2155]  = 1;
  ram[2156]  = 1;
  ram[2157]  = 1;
  ram[2158]  = 1;
  ram[2159]  = 1;
  ram[2160]  = 1;
  ram[2161]  = 1;
  ram[2162]  = 1;
  ram[2163]  = 1;
  ram[2164]  = 1;
  ram[2165]  = 1;
  ram[2166]  = 1;
  ram[2167]  = 1;
  ram[2168]  = 1;
  ram[2169]  = 1;
  ram[2170]  = 1;
  ram[2171]  = 1;
  ram[2172]  = 1;
  ram[2173]  = 1;
  ram[2174]  = 1;
  ram[2175]  = 1;
  ram[2176]  = 1;
  ram[2177]  = 1;
  ram[2178]  = 1;
  ram[2179]  = 1;
  ram[2180]  = 1;
  ram[2181]  = 1;
  ram[2182]  = 1;
  ram[2183]  = 1;
  ram[2184]  = 1;
  ram[2185]  = 1;
  ram[2186]  = 1;
  ram[2187]  = 1;
  ram[2188]  = 1;
  ram[2189]  = 1;
  ram[2190]  = 1;
  ram[2191]  = 1;
  ram[2192]  = 1;
  ram[2193]  = 1;
  ram[2194]  = 1;
  ram[2195]  = 1;
  ram[2196]  = 1;
  ram[2197]  = 1;
  ram[2198]  = 1;
  ram[2199]  = 1;
  ram[2200]  = 1;
  ram[2201]  = 1;
  ram[2202]  = 1;
  ram[2203]  = 1;
  ram[2204]  = 1;
  ram[2205]  = 1;
  ram[2206]  = 1;
  ram[2207]  = 1;
  ram[2208]  = 1;
  ram[2209]  = 1;
  ram[2210]  = 1;
  ram[2211]  = 1;
  ram[2212]  = 1;
  ram[2213]  = 1;
  ram[2214]  = 1;
  ram[2215]  = 1;
  ram[2216]  = 1;
  ram[2217]  = 1;
  ram[2218]  = 1;
  ram[2219]  = 1;
  ram[2220]  = 1;
  ram[2221]  = 1;
  ram[2222]  = 1;
  ram[2223]  = 1;
  ram[2224]  = 1;
  ram[2225]  = 1;
  ram[2226]  = 1;
  ram[2227]  = 1;
  ram[2228]  = 1;
  ram[2229]  = 1;
  ram[2230]  = 1;
  ram[2231]  = 1;
  ram[2232]  = 1;
  ram[2233]  = 1;
  ram[2234]  = 1;
  ram[2235]  = 1;
  ram[2236]  = 1;
  ram[2237]  = 1;
  ram[2238]  = 1;
  ram[2239]  = 1;
  ram[2240]  = 1;
  ram[2241]  = 1;
  ram[2242]  = 1;
  ram[2243]  = 1;
  ram[2244]  = 1;
  ram[2245]  = 1;
  ram[2246]  = 1;
  ram[2247]  = 1;
  ram[2248]  = 1;
  ram[2249]  = 1;
  ram[2250]  = 1;
  ram[2251]  = 1;
  ram[2252]  = 1;
  ram[2253]  = 1;
  ram[2254]  = 1;
  ram[2255]  = 1;
  ram[2256]  = 1;
  ram[2257]  = 1;
  ram[2258]  = 1;
  ram[2259]  = 1;
  ram[2260]  = 1;
  ram[2261]  = 1;
  ram[2262]  = 1;
  ram[2263]  = 1;
  ram[2264]  = 1;
  ram[2265]  = 1;
  ram[2266]  = 1;
  ram[2267]  = 1;
  ram[2268]  = 1;
  ram[2269]  = 1;
  ram[2270]  = 1;
  ram[2271]  = 1;
  ram[2272]  = 1;
  ram[2273]  = 1;
  ram[2274]  = 1;
  ram[2275]  = 1;
  ram[2276]  = 1;
  ram[2277]  = 1;
  ram[2278]  = 1;
  ram[2279]  = 1;
  ram[2280]  = 1;
  ram[2281]  = 1;
  ram[2282]  = 1;
  ram[2283]  = 1;
  ram[2284]  = 1;
  ram[2285]  = 1;
  ram[2286]  = 1;
  ram[2287]  = 1;
  ram[2288]  = 1;
  ram[2289]  = 1;
  ram[2290]  = 1;
  ram[2291]  = 1;
  ram[2292]  = 1;
  ram[2293]  = 1;
  ram[2294]  = 1;
  ram[2295]  = 1;
  ram[2296]  = 1;
  ram[2297]  = 1;
  ram[2298]  = 1;
  ram[2299]  = 1;
  ram[2300]  = 1;
  ram[2301]  = 1;
  ram[2302]  = 1;
  ram[2303]  = 1;
  ram[2304]  = 1;
  ram[2305]  = 1;
  ram[2306]  = 1;
  ram[2307]  = 1;
  ram[2308]  = 1;
  ram[2309]  = 1;
  ram[2310]  = 1;
  ram[2311]  = 1;
  ram[2312]  = 1;
  ram[2313]  = 1;
  ram[2314]  = 1;
  ram[2315]  = 1;
  ram[2316]  = 1;
  ram[2317]  = 1;
  ram[2318]  = 1;
  ram[2319]  = 1;
  ram[2320]  = 1;
  ram[2321]  = 1;
  ram[2322]  = 1;
  ram[2323]  = 1;
  ram[2324]  = 1;
  ram[2325]  = 1;
  ram[2326]  = 1;
  ram[2327]  = 1;
  ram[2328]  = 1;
  ram[2329]  = 1;
  ram[2330]  = 1;
  ram[2331]  = 1;
  ram[2332]  = 1;
  ram[2333]  = 1;
  ram[2334]  = 1;
  ram[2335]  = 1;
  ram[2336]  = 1;
  ram[2337]  = 1;
  ram[2338]  = 1;
  ram[2339]  = 1;
  ram[2340]  = 1;
  ram[2341]  = 1;
  ram[2342]  = 1;
  ram[2343]  = 1;
  ram[2344]  = 1;
  ram[2345]  = 1;
  ram[2346]  = 1;
  ram[2347]  = 1;
  ram[2348]  = 1;
  ram[2349]  = 1;
  ram[2350]  = 1;
  ram[2351]  = 1;
  ram[2352]  = 1;
  ram[2353]  = 1;
  ram[2354]  = 1;
  ram[2355]  = 1;
  ram[2356]  = 1;
  ram[2357]  = 1;
  ram[2358]  = 1;
  ram[2359]  = 1;
  ram[2360]  = 1;
  ram[2361]  = 1;
  ram[2362]  = 1;
  ram[2363]  = 1;
  ram[2364]  = 1;
  ram[2365]  = 1;
  ram[2366]  = 1;
  ram[2367]  = 1;
  ram[2368]  = 1;
  ram[2369]  = 1;
  ram[2370]  = 1;
  ram[2371]  = 1;
  ram[2372]  = 1;
  ram[2373]  = 1;
  ram[2374]  = 1;
  ram[2375]  = 1;
  ram[2376]  = 1;
  ram[2377]  = 1;
  ram[2378]  = 1;
  ram[2379]  = 1;
  ram[2380]  = 1;
  ram[2381]  = 1;
  ram[2382]  = 1;
  ram[2383]  = 1;
  ram[2384]  = 1;
  ram[2385]  = 1;
  ram[2386]  = 1;
  ram[2387]  = 1;
  ram[2388]  = 1;
  ram[2389]  = 1;
  ram[2390]  = 1;
  ram[2391]  = 1;
  ram[2392]  = 1;
  ram[2393]  = 1;
  ram[2394]  = 1;
  ram[2395]  = 1;
  ram[2396]  = 1;
  ram[2397]  = 1;
  ram[2398]  = 1;
  ram[2399]  = 1;
  ram[2400]  = 1;
  ram[2401]  = 1;
  ram[2402]  = 1;
  ram[2403]  = 1;
  ram[2404]  = 1;
  ram[2405]  = 1;
  ram[2406]  = 1;
  ram[2407]  = 1;
  ram[2408]  = 1;
  ram[2409]  = 1;
  ram[2410]  = 1;
  ram[2411]  = 1;
  ram[2412]  = 1;
  ram[2413]  = 1;
  ram[2414]  = 1;
  ram[2415]  = 1;
  ram[2416]  = 1;
  ram[2417]  = 1;
  ram[2418]  = 1;
  ram[2419]  = 1;
  ram[2420]  = 1;
  ram[2421]  = 1;
  ram[2422]  = 1;
  ram[2423]  = 1;
  ram[2424]  = 1;
  ram[2425]  = 1;
  ram[2426]  = 1;
  ram[2427]  = 1;
  ram[2428]  = 1;
  ram[2429]  = 1;
  ram[2430]  = 1;
  ram[2431]  = 1;
  ram[2432]  = 1;
  ram[2433]  = 1;
  ram[2434]  = 1;
  ram[2435]  = 1;
  ram[2436]  = 1;
  ram[2437]  = 1;
  ram[2438]  = 1;
  ram[2439]  = 1;
  ram[2440]  = 1;
  ram[2441]  = 1;
  ram[2442]  = 1;
  ram[2443]  = 1;
  ram[2444]  = 1;
  ram[2445]  = 1;
  ram[2446]  = 1;
  ram[2447]  = 1;
  ram[2448]  = 1;
  ram[2449]  = 1;
  ram[2450]  = 1;
  ram[2451]  = 1;
  ram[2452]  = 1;
  ram[2453]  = 1;
  ram[2454]  = 1;
  ram[2455]  = 1;
  ram[2456]  = 1;
  ram[2457]  = 1;
  ram[2458]  = 1;
  ram[2459]  = 1;
  ram[2460]  = 1;
  ram[2461]  = 1;
  ram[2462]  = 1;
  ram[2463]  = 1;
  ram[2464]  = 1;
  ram[2465]  = 1;
  ram[2466]  = 1;
  ram[2467]  = 1;
  ram[2468]  = 1;
  ram[2469]  = 1;
  ram[2470]  = 1;
  ram[2471]  = 1;
  ram[2472]  = 1;
  ram[2473]  = 1;
  ram[2474]  = 1;
  ram[2475]  = 1;
  ram[2476]  = 1;
  ram[2477]  = 1;
  ram[2478]  = 1;
  ram[2479]  = 1;
  ram[2480]  = 1;
  ram[2481]  = 1;
  ram[2482]  = 1;
  ram[2483]  = 1;
  ram[2484]  = 1;
  ram[2485]  = 1;
  ram[2486]  = 1;
  ram[2487]  = 1;
  ram[2488]  = 1;
  ram[2489]  = 1;
  ram[2490]  = 1;
  ram[2491]  = 1;
  ram[2492]  = 1;
  ram[2493]  = 1;
  ram[2494]  = 1;
  ram[2495]  = 1;
  ram[2496]  = 1;
  ram[2497]  = 1;
  ram[2498]  = 1;
  ram[2499]  = 1;
  ram[2500]  = 1;
  ram[2501]  = 1;
  ram[2502]  = 1;
  ram[2503]  = 1;
  ram[2504]  = 1;
  ram[2505]  = 1;
  ram[2506]  = 1;
  ram[2507]  = 1;
  ram[2508]  = 1;
  ram[2509]  = 1;
  ram[2510]  = 1;
  ram[2511]  = 1;
  ram[2512]  = 1;
  ram[2513]  = 1;
  ram[2514]  = 1;
  ram[2515]  = 1;
  ram[2516]  = 1;
  ram[2517]  = 1;
  ram[2518]  = 1;
  ram[2519]  = 1;
  ram[2520]  = 1;
  ram[2521]  = 1;
  ram[2522]  = 1;
  ram[2523]  = 1;
  ram[2524]  = 1;
  ram[2525]  = 1;
  ram[2526]  = 1;
  ram[2527]  = 1;
  ram[2528]  = 1;
  ram[2529]  = 1;
  ram[2530]  = 1;
  ram[2531]  = 1;
  ram[2532]  = 1;
  ram[2533]  = 1;
  ram[2534]  = 1;
  ram[2535]  = 1;
  ram[2536]  = 1;
  ram[2537]  = 1;
  ram[2538]  = 1;
  ram[2539]  = 1;
  ram[2540]  = 1;
  ram[2541]  = 1;
  ram[2542]  = 1;
  ram[2543]  = 1;
  ram[2544]  = 1;
  ram[2545]  = 1;
  ram[2546]  = 1;
  ram[2547]  = 1;
  ram[2548]  = 1;
  ram[2549]  = 1;
  ram[2550]  = 1;
  ram[2551]  = 1;
  ram[2552]  = 1;
  ram[2553]  = 1;
  ram[2554]  = 1;
  ram[2555]  = 1;
  ram[2556]  = 1;
  ram[2557]  = 1;
  ram[2558]  = 1;
  ram[2559]  = 1;
  ram[2560]  = 1;
  ram[2561]  = 1;
  ram[2562]  = 1;
  ram[2563]  = 1;
  ram[2564]  = 1;
  ram[2565]  = 1;
  ram[2566]  = 1;
  ram[2567]  = 1;
  ram[2568]  = 1;
  ram[2569]  = 1;
  ram[2570]  = 1;
  ram[2571]  = 1;
  ram[2572]  = 1;
  ram[2573]  = 1;
  ram[2574]  = 1;
  ram[2575]  = 1;
  ram[2576]  = 1;
  ram[2577]  = 1;
  ram[2578]  = 1;
  ram[2579]  = 1;
  ram[2580]  = 1;
  ram[2581]  = 1;
  ram[2582]  = 1;
  ram[2583]  = 1;
  ram[2584]  = 1;
  ram[2585]  = 1;
  ram[2586]  = 1;
  ram[2587]  = 1;
  ram[2588]  = 1;
  ram[2589]  = 1;
  ram[2590]  = 1;
  ram[2591]  = 1;
  ram[2592]  = 1;
  ram[2593]  = 1;
  ram[2594]  = 1;
  ram[2595]  = 1;
  ram[2596]  = 1;
  ram[2597]  = 1;
  ram[2598]  = 1;
  ram[2599]  = 1;
  ram[2600]  = 1;
  ram[2601]  = 1;
  ram[2602]  = 1;
  ram[2603]  = 1;
  ram[2604]  = 1;
  ram[2605]  = 1;
  ram[2606]  = 1;
  ram[2607]  = 1;
  ram[2608]  = 1;
  ram[2609]  = 1;
  ram[2610]  = 1;
  ram[2611]  = 1;
  ram[2612]  = 1;
  ram[2613]  = 1;
  ram[2614]  = 1;
  ram[2615]  = 1;
  ram[2616]  = 1;
  ram[2617]  = 1;
  ram[2618]  = 1;
  ram[2619]  = 1;
  ram[2620]  = 1;
  ram[2621]  = 1;
  ram[2622]  = 1;
  ram[2623]  = 1;
  ram[2624]  = 1;
  ram[2625]  = 1;
  ram[2626]  = 1;
  ram[2627]  = 1;
  ram[2628]  = 1;
  ram[2629]  = 1;
  ram[2630]  = 1;
  ram[2631]  = 1;
  ram[2632]  = 1;
  ram[2633]  = 1;
  ram[2634]  = 1;
  ram[2635]  = 1;
  ram[2636]  = 1;
  ram[2637]  = 1;
  ram[2638]  = 1;
  ram[2639]  = 1;
  ram[2640]  = 1;
  ram[2641]  = 1;
  ram[2642]  = 1;
  ram[2643]  = 1;
  ram[2644]  = 1;
  ram[2645]  = 1;
  ram[2646]  = 1;
  ram[2647]  = 1;
  ram[2648]  = 1;
  ram[2649]  = 1;
  ram[2650]  = 1;
  ram[2651]  = 1;
  ram[2652]  = 1;
  ram[2653]  = 1;
  ram[2654]  = 1;
  ram[2655]  = 1;
  ram[2656]  = 1;
  ram[2657]  = 1;
  ram[2658]  = 1;
  ram[2659]  = 1;
  ram[2660]  = 1;
  ram[2661]  = 1;
  ram[2662]  = 1;
  ram[2663]  = 1;
  ram[2664]  = 1;
  ram[2665]  = 1;
  ram[2666]  = 1;
  ram[2667]  = 1;
  ram[2668]  = 1;
  ram[2669]  = 1;
  ram[2670]  = 1;
  ram[2671]  = 1;
  ram[2672]  = 1;
  ram[2673]  = 1;
  ram[2674]  = 1;
  ram[2675]  = 1;
  ram[2676]  = 1;
  ram[2677]  = 1;
  ram[2678]  = 1;
  ram[2679]  = 1;
  ram[2680]  = 1;
  ram[2681]  = 1;
  ram[2682]  = 1;
  ram[2683]  = 1;
  ram[2684]  = 1;
  ram[2685]  = 1;
  ram[2686]  = 1;
  ram[2687]  = 1;
  ram[2688]  = 1;
  ram[2689]  = 1;
  ram[2690]  = 1;
  ram[2691]  = 1;
  ram[2692]  = 1;
  ram[2693]  = 1;
  ram[2694]  = 1;
  ram[2695]  = 1;
  ram[2696]  = 1;
  ram[2697]  = 1;
  ram[2698]  = 1;
  ram[2699]  = 1;
  ram[2700]  = 1;
  ram[2701]  = 1;
  ram[2702]  = 1;
  ram[2703]  = 1;
  ram[2704]  = 1;
  ram[2705]  = 1;
  ram[2706]  = 1;
  ram[2707]  = 1;
  ram[2708]  = 1;
  ram[2709]  = 1;
  ram[2710]  = 1;
  ram[2711]  = 1;
  ram[2712]  = 1;
  ram[2713]  = 1;
  ram[2714]  = 1;
  ram[2715]  = 1;
  ram[2716]  = 1;
  ram[2717]  = 1;
  ram[2718]  = 1;
  ram[2719]  = 1;
  ram[2720]  = 1;
  ram[2721]  = 1;
  ram[2722]  = 1;
  ram[2723]  = 1;
  ram[2724]  = 1;
  ram[2725]  = 1;
  ram[2726]  = 1;
  ram[2727]  = 1;
  ram[2728]  = 1;
  ram[2729]  = 1;
  ram[2730]  = 1;
  ram[2731]  = 1;
  ram[2732]  = 1;
  ram[2733]  = 1;
  ram[2734]  = 1;
  ram[2735]  = 1;
  ram[2736]  = 1;
  ram[2737]  = 1;
  ram[2738]  = 1;
  ram[2739]  = 1;
  ram[2740]  = 1;
  ram[2741]  = 1;
  ram[2742]  = 1;
  ram[2743]  = 1;
  ram[2744]  = 1;
  ram[2745]  = 1;
  ram[2746]  = 1;
  ram[2747]  = 1;
  ram[2748]  = 1;
  ram[2749]  = 1;
  ram[2750]  = 1;
  ram[2751]  = 1;
  ram[2752]  = 1;
  ram[2753]  = 1;
  ram[2754]  = 1;
  ram[2755]  = 1;
  ram[2756]  = 1;
  ram[2757]  = 1;
  ram[2758]  = 1;
  ram[2759]  = 1;
  ram[2760]  = 1;
  ram[2761]  = 1;
  ram[2762]  = 1;
  ram[2763]  = 1;
  ram[2764]  = 1;
  ram[2765]  = 1;
  ram[2766]  = 1;
  ram[2767]  = 1;
  ram[2768]  = 1;
  ram[2769]  = 1;
  ram[2770]  = 1;
  ram[2771]  = 1;
  ram[2772]  = 1;
  ram[2773]  = 1;
  ram[2774]  = 1;
  ram[2775]  = 1;
  ram[2776]  = 1;
  ram[2777]  = 1;
  ram[2778]  = 1;
  ram[2779]  = 1;
  ram[2780]  = 1;
  ram[2781]  = 1;
  ram[2782]  = 1;
  ram[2783]  = 1;
  ram[2784]  = 1;
  ram[2785]  = 1;
  ram[2786]  = 1;
  ram[2787]  = 1;
  ram[2788]  = 1;
  ram[2789]  = 1;
  ram[2790]  = 1;
  ram[2791]  = 1;
  ram[2792]  = 1;
  ram[2793]  = 1;
  ram[2794]  = 1;
  ram[2795]  = 1;
  ram[2796]  = 1;
  ram[2797]  = 1;
  ram[2798]  = 1;
  ram[2799]  = 1;
  ram[2800]  = 1;
  ram[2801]  = 1;
  ram[2802]  = 1;
  ram[2803]  = 1;
  ram[2804]  = 1;
  ram[2805]  = 1;
  ram[2806]  = 1;
  ram[2807]  = 1;
  ram[2808]  = 1;
  ram[2809]  = 1;
  ram[2810]  = 1;
  ram[2811]  = 1;
  ram[2812]  = 1;
  ram[2813]  = 1;
  ram[2814]  = 1;
  ram[2815]  = 1;
  ram[2816]  = 1;
  ram[2817]  = 1;
  ram[2818]  = 1;
  ram[2819]  = 1;
  ram[2820]  = 1;
  ram[2821]  = 1;
  ram[2822]  = 1;
  ram[2823]  = 1;
  ram[2824]  = 1;
  ram[2825]  = 1;
  ram[2826]  = 1;
  ram[2827]  = 1;
  ram[2828]  = 1;
  ram[2829]  = 1;
  ram[2830]  = 1;
  ram[2831]  = 1;
  ram[2832]  = 1;
  ram[2833]  = 1;
  ram[2834]  = 1;
  ram[2835]  = 1;
  ram[2836]  = 1;
  ram[2837]  = 1;
  ram[2838]  = 1;
  ram[2839]  = 1;
  ram[2840]  = 1;
  ram[2841]  = 1;
  ram[2842]  = 1;
  ram[2843]  = 1;
  ram[2844]  = 1;
  ram[2845]  = 1;
  ram[2846]  = 1;
  ram[2847]  = 1;
  ram[2848]  = 1;
  ram[2849]  = 1;
  ram[2850]  = 1;
  ram[2851]  = 1;
  ram[2852]  = 1;
  ram[2853]  = 1;
  ram[2854]  = 1;
  ram[2855]  = 1;
  ram[2856]  = 1;
  ram[2857]  = 1;
  ram[2858]  = 1;
  ram[2859]  = 1;
  ram[2860]  = 1;
  ram[2861]  = 1;
  ram[2862]  = 1;
  ram[2863]  = 1;
  ram[2864]  = 1;
  ram[2865]  = 1;
  ram[2866]  = 1;
  ram[2867]  = 1;
  ram[2868]  = 1;
  ram[2869]  = 1;
  ram[2870]  = 1;
  ram[2871]  = 1;
  ram[2872]  = 1;
  ram[2873]  = 1;
  ram[2874]  = 1;
  ram[2875]  = 1;
  ram[2876]  = 1;
  ram[2877]  = 1;
  ram[2878]  = 1;
  ram[2879]  = 1;
  ram[2880]  = 1;
  ram[2881]  = 1;
  ram[2882]  = 1;
  ram[2883]  = 1;
  ram[2884]  = 1;
  ram[2885]  = 1;
  ram[2886]  = 1;
  ram[2887]  = 1;
  ram[2888]  = 1;
  ram[2889]  = 1;
  ram[2890]  = 1;
  ram[2891]  = 1;
  ram[2892]  = 1;
  ram[2893]  = 1;
  ram[2894]  = 1;
  ram[2895]  = 1;
  ram[2896]  = 1;
  ram[2897]  = 1;
  ram[2898]  = 1;
  ram[2899]  = 1;
  ram[2900]  = 1;
  ram[2901]  = 1;
  ram[2902]  = 1;
  ram[2903]  = 1;
  ram[2904]  = 1;
  ram[2905]  = 1;
  ram[2906]  = 1;
  ram[2907]  = 1;
  ram[2908]  = 1;
  ram[2909]  = 1;
  ram[2910]  = 1;
  ram[2911]  = 1;
  ram[2912]  = 1;
  ram[2913]  = 1;
  ram[2914]  = 1;
  ram[2915]  = 1;
  ram[2916]  = 1;
  ram[2917]  = 1;
  ram[2918]  = 1;
  ram[2919]  = 1;
  ram[2920]  = 1;
  ram[2921]  = 1;
  ram[2922]  = 1;
  ram[2923]  = 1;
  ram[2924]  = 1;
  ram[2925]  = 1;
  ram[2926]  = 1;
  ram[2927]  = 1;
  ram[2928]  = 1;
  ram[2929]  = 1;
  ram[2930]  = 1;
  ram[2931]  = 1;
  ram[2932]  = 1;
  ram[2933]  = 1;
  ram[2934]  = 1;
  ram[2935]  = 1;
  ram[2936]  = 1;
  ram[2937]  = 1;
  ram[2938]  = 1;
  ram[2939]  = 1;
  ram[2940]  = 1;
  ram[2941]  = 1;
  ram[2942]  = 1;
  ram[2943]  = 1;
  ram[2944]  = 1;
  ram[2945]  = 1;
  ram[2946]  = 1;
  ram[2947]  = 1;
  ram[2948]  = 1;
  ram[2949]  = 1;
  ram[2950]  = 1;
  ram[2951]  = 1;
  ram[2952]  = 1;
  ram[2953]  = 1;
  ram[2954]  = 1;
  ram[2955]  = 1;
  ram[2956]  = 1;
  ram[2957]  = 1;
  ram[2958]  = 1;
  ram[2959]  = 1;
  ram[2960]  = 1;
  ram[2961]  = 1;
  ram[2962]  = 1;
  ram[2963]  = 1;
  ram[2964]  = 1;
  ram[2965]  = 1;
  ram[2966]  = 1;
  ram[2967]  = 1;
  ram[2968]  = 1;
  ram[2969]  = 1;
  ram[2970]  = 1;
  ram[2971]  = 1;
  ram[2972]  = 1;
  ram[2973]  = 1;
  ram[2974]  = 1;
  ram[2975]  = 1;
  ram[2976]  = 1;
  ram[2977]  = 1;
  ram[2978]  = 1;
  ram[2979]  = 1;
  ram[2980]  = 1;
  ram[2981]  = 1;
  ram[2982]  = 1;
  ram[2983]  = 1;
  ram[2984]  = 1;
  ram[2985]  = 1;
  ram[2986]  = 1;
  ram[2987]  = 1;
  ram[2988]  = 1;
  ram[2989]  = 1;
  ram[2990]  = 1;
  ram[2991]  = 1;
  ram[2992]  = 1;
  ram[2993]  = 1;
  ram[2994]  = 1;
  ram[2995]  = 1;
  ram[2996]  = 1;
  ram[2997]  = 1;
  ram[2998]  = 1;
  ram[2999]  = 1;
  ram[3000]  = 1;
  ram[3001]  = 1;
  ram[3002]  = 1;
  ram[3003]  = 1;
  ram[3004]  = 1;
  ram[3005]  = 1;
  ram[3006]  = 1;
  ram[3007]  = 1;
  ram[3008]  = 1;
  ram[3009]  = 1;
  ram[3010]  = 1;
  ram[3011]  = 1;
  ram[3012]  = 1;
  ram[3013]  = 1;
  ram[3014]  = 1;
  ram[3015]  = 1;
  ram[3016]  = 1;
  ram[3017]  = 1;
  ram[3018]  = 1;
  ram[3019]  = 1;
  ram[3020]  = 1;
  ram[3021]  = 1;
  ram[3022]  = 1;
  ram[3023]  = 1;
  ram[3024]  = 1;
  ram[3025]  = 1;
  ram[3026]  = 1;
  ram[3027]  = 1;
  ram[3028]  = 1;
  ram[3029]  = 1;
  ram[3030]  = 1;
  ram[3031]  = 1;
  ram[3032]  = 1;
  ram[3033]  = 1;
  ram[3034]  = 1;
  ram[3035]  = 1;
  ram[3036]  = 1;
  ram[3037]  = 1;
  ram[3038]  = 1;
  ram[3039]  = 1;
  ram[3040]  = 1;
  ram[3041]  = 1;
  ram[3042]  = 1;
  ram[3043]  = 1;
  ram[3044]  = 1;
  ram[3045]  = 1;
  ram[3046]  = 1;
  ram[3047]  = 1;
  ram[3048]  = 1;
  ram[3049]  = 1;
  ram[3050]  = 1;
  ram[3051]  = 1;
  ram[3052]  = 1;
  ram[3053]  = 1;
  ram[3054]  = 1;
  ram[3055]  = 1;
  ram[3056]  = 1;
  ram[3057]  = 1;
  ram[3058]  = 1;
  ram[3059]  = 1;
  ram[3060]  = 1;
  ram[3061]  = 1;
  ram[3062]  = 1;
  ram[3063]  = 1;
  ram[3064]  = 1;
  ram[3065]  = 1;
  ram[3066]  = 1;
  ram[3067]  = 1;
  ram[3068]  = 1;
  ram[3069]  = 1;
  ram[3070]  = 1;
  ram[3071]  = 1;
  ram[3072]  = 1;
  ram[3073]  = 1;
  ram[3074]  = 1;
  ram[3075]  = 1;
  ram[3076]  = 1;
  ram[3077]  = 1;
  ram[3078]  = 1;
  ram[3079]  = 1;
  ram[3080]  = 1;
  ram[3081]  = 1;
  ram[3082]  = 1;
  ram[3083]  = 1;
  ram[3084]  = 1;
  ram[3085]  = 1;
  ram[3086]  = 1;
  ram[3087]  = 1;
  ram[3088]  = 1;
  ram[3089]  = 1;
  ram[3090]  = 1;
  ram[3091]  = 1;
  ram[3092]  = 1;
  ram[3093]  = 1;
  ram[3094]  = 1;
  ram[3095]  = 1;
  ram[3096]  = 1;
  ram[3097]  = 1;
  ram[3098]  = 1;
  ram[3099]  = 1;
  ram[3100]  = 1;
  ram[3101]  = 1;
  ram[3102]  = 1;
  ram[3103]  = 1;
  ram[3104]  = 1;
  ram[3105]  = 1;
  ram[3106]  = 1;
  ram[3107]  = 1;
  ram[3108]  = 1;
  ram[3109]  = 1;
  ram[3110]  = 1;
  ram[3111]  = 1;
  ram[3112]  = 1;
  ram[3113]  = 1;
  ram[3114]  = 1;
  ram[3115]  = 1;
  ram[3116]  = 1;
  ram[3117]  = 1;
  ram[3118]  = 1;
  ram[3119]  = 1;
  ram[3120]  = 1;
  ram[3121]  = 1;
  ram[3122]  = 1;
  ram[3123]  = 1;
  ram[3124]  = 1;
  ram[3125]  = 1;
  ram[3126]  = 1;
  ram[3127]  = 1;
  ram[3128]  = 1;
  ram[3129]  = 1;
  ram[3130]  = 1;
  ram[3131]  = 1;
  ram[3132]  = 1;
  ram[3133]  = 1;
  ram[3134]  = 1;
  ram[3135]  = 1;
  ram[3136]  = 1;
  ram[3137]  = 1;
  ram[3138]  = 1;
  ram[3139]  = 1;
  ram[3140]  = 1;
  ram[3141]  = 1;
  ram[3142]  = 1;
  ram[3143]  = 1;
  ram[3144]  = 1;
  ram[3145]  = 1;
  ram[3146]  = 1;
  ram[3147]  = 1;
  ram[3148]  = 1;
  ram[3149]  = 1;
  ram[3150]  = 1;
  ram[3151]  = 1;
  ram[3152]  = 1;
  ram[3153]  = 1;
  ram[3154]  = 1;
  ram[3155]  = 1;
  ram[3156]  = 1;
  ram[3157]  = 1;
  ram[3158]  = 1;
  ram[3159]  = 1;
  ram[3160]  = 1;
  ram[3161]  = 1;
  ram[3162]  = 1;
  ram[3163]  = 1;
  ram[3164]  = 1;
  ram[3165]  = 1;
  ram[3166]  = 1;
  ram[3167]  = 1;
  ram[3168]  = 1;
  ram[3169]  = 1;
  ram[3170]  = 1;
  ram[3171]  = 1;
  ram[3172]  = 1;
  ram[3173]  = 1;
  ram[3174]  = 1;
  ram[3175]  = 1;
  ram[3176]  = 1;
  ram[3177]  = 1;
  ram[3178]  = 1;
  ram[3179]  = 1;
  ram[3180]  = 1;
  ram[3181]  = 1;
  ram[3182]  = 1;
  ram[3183]  = 1;
  ram[3184]  = 1;
  ram[3185]  = 1;
  ram[3186]  = 1;
  ram[3187]  = 1;
  ram[3188]  = 1;
  ram[3189]  = 1;
  ram[3190]  = 1;
  ram[3191]  = 1;
  ram[3192]  = 1;
  ram[3193]  = 1;
  ram[3194]  = 1;
  ram[3195]  = 1;
  ram[3196]  = 1;
  ram[3197]  = 1;
  ram[3198]  = 1;
  ram[3199]  = 1;
  ram[3200]  = 1;
  ram[3201]  = 1;
  ram[3202]  = 1;
  ram[3203]  = 1;
  ram[3204]  = 1;
  ram[3205]  = 1;
  ram[3206]  = 1;
  ram[3207]  = 1;
  ram[3208]  = 1;
  ram[3209]  = 1;
  ram[3210]  = 1;
  ram[3211]  = 1;
  ram[3212]  = 1;
  ram[3213]  = 1;
  ram[3214]  = 1;
  ram[3215]  = 1;
  ram[3216]  = 1;
  ram[3217]  = 1;
  ram[3218]  = 1;
  ram[3219]  = 1;
  ram[3220]  = 1;
  ram[3221]  = 1;
  ram[3222]  = 1;
  ram[3223]  = 1;
  ram[3224]  = 1;
  ram[3225]  = 1;
  ram[3226]  = 1;
  ram[3227]  = 1;
  ram[3228]  = 1;
  ram[3229]  = 1;
  ram[3230]  = 1;
  ram[3231]  = 1;
  ram[3232]  = 1;
  ram[3233]  = 1;
  ram[3234]  = 1;
  ram[3235]  = 1;
  ram[3236]  = 1;
  ram[3237]  = 1;
  ram[3238]  = 1;
  ram[3239]  = 1;
  ram[3240]  = 1;
  ram[3241]  = 1;
  ram[3242]  = 1;
  ram[3243]  = 1;
  ram[3244]  = 1;
  ram[3245]  = 1;
  ram[3246]  = 1;
  ram[3247]  = 1;
  ram[3248]  = 1;
  ram[3249]  = 1;
  ram[3250]  = 1;
  ram[3251]  = 1;
  ram[3252]  = 1;
  ram[3253]  = 1;
  ram[3254]  = 1;
  ram[3255]  = 1;
  ram[3256]  = 1;
  ram[3257]  = 1;
  ram[3258]  = 1;
  ram[3259]  = 1;
  ram[3260]  = 1;
  ram[3261]  = 1;
  ram[3262]  = 1;
  ram[3263]  = 1;
  ram[3264]  = 1;
  ram[3265]  = 1;
  ram[3266]  = 1;
  ram[3267]  = 1;
  ram[3268]  = 1;
  ram[3269]  = 1;
  ram[3270]  = 1;
  ram[3271]  = 1;
  ram[3272]  = 1;
  ram[3273]  = 1;
  ram[3274]  = 1;
  ram[3275]  = 1;
  ram[3276]  = 1;
  ram[3277]  = 1;
  ram[3278]  = 1;
  ram[3279]  = 1;
  ram[3280]  = 1;
  ram[3281]  = 1;
  ram[3282]  = 1;
  ram[3283]  = 1;
  ram[3284]  = 1;
  ram[3285]  = 1;
  ram[3286]  = 1;
  ram[3287]  = 1;
  ram[3288]  = 1;
  ram[3289]  = 1;
  ram[3290]  = 1;
  ram[3291]  = 1;
  ram[3292]  = 1;
  ram[3293]  = 1;
  ram[3294]  = 1;
  ram[3295]  = 1;
  ram[3296]  = 1;
  ram[3297]  = 1;
  ram[3298]  = 1;
  ram[3299]  = 1;
  ram[3300]  = 1;
  ram[3301]  = 1;
  ram[3302]  = 1;
  ram[3303]  = 1;
  ram[3304]  = 1;
  ram[3305]  = 1;
  ram[3306]  = 1;
  ram[3307]  = 1;
  ram[3308]  = 1;
  ram[3309]  = 1;
  ram[3310]  = 1;
  ram[3311]  = 1;
  ram[3312]  = 1;
  ram[3313]  = 1;
  ram[3314]  = 1;
  ram[3315]  = 1;
  ram[3316]  = 1;
  ram[3317]  = 1;
  ram[3318]  = 1;
  ram[3319]  = 1;
  ram[3320]  = 1;
  ram[3321]  = 1;
  ram[3322]  = 1;
  ram[3323]  = 1;
  ram[3324]  = 1;
  ram[3325]  = 1;
  ram[3326]  = 1;
  ram[3327]  = 1;
  ram[3328]  = 1;
  ram[3329]  = 1;
  ram[3330]  = 1;
  ram[3331]  = 1;
  ram[3332]  = 1;
  ram[3333]  = 1;
  ram[3334]  = 1;
  ram[3335]  = 1;
  ram[3336]  = 1;
  ram[3337]  = 1;
  ram[3338]  = 1;
  ram[3339]  = 1;
  ram[3340]  = 1;
  ram[3341]  = 1;
  ram[3342]  = 1;
  ram[3343]  = 1;
  ram[3344]  = 1;
  ram[3345]  = 1;
  ram[3346]  = 1;
  ram[3347]  = 1;
  ram[3348]  = 1;
  ram[3349]  = 1;
  ram[3350]  = 1;
  ram[3351]  = 1;
  ram[3352]  = 1;
  ram[3353]  = 1;
  ram[3354]  = 1;
  ram[3355]  = 1;
  ram[3356]  = 1;
  ram[3357]  = 1;
  ram[3358]  = 1;
  ram[3359]  = 1;
  ram[3360]  = 1;
  ram[3361]  = 1;
  ram[3362]  = 1;
  ram[3363]  = 1;
  ram[3364]  = 1;
  ram[3365]  = 1;
  ram[3366]  = 1;
  ram[3367]  = 1;
  ram[3368]  = 1;
  ram[3369]  = 1;
  ram[3370]  = 1;
  ram[3371]  = 1;
  ram[3372]  = 1;
  ram[3373]  = 1;
  ram[3374]  = 1;
  ram[3375]  = 1;
  ram[3376]  = 1;
  ram[3377]  = 1;
  ram[3378]  = 1;
  ram[3379]  = 1;
  ram[3380]  = 1;
  ram[3381]  = 1;
  ram[3382]  = 1;
  ram[3383]  = 1;
  ram[3384]  = 1;
  ram[3385]  = 1;
  ram[3386]  = 1;
  ram[3387]  = 1;
  ram[3388]  = 1;
  ram[3389]  = 1;
  ram[3390]  = 1;
  ram[3391]  = 1;
  ram[3392]  = 1;
  ram[3393]  = 1;
  ram[3394]  = 1;
  ram[3395]  = 1;
  ram[3396]  = 1;
  ram[3397]  = 1;
  ram[3398]  = 1;
  ram[3399]  = 1;
  ram[3400]  = 1;
  ram[3401]  = 1;
  ram[3402]  = 1;
  ram[3403]  = 1;
  ram[3404]  = 1;
  ram[3405]  = 1;
  ram[3406]  = 1;
  ram[3407]  = 1;
  ram[3408]  = 1;
  ram[3409]  = 1;
  ram[3410]  = 1;
  ram[3411]  = 1;
  ram[3412]  = 1;
  ram[3413]  = 1;
  ram[3414]  = 1;
  ram[3415]  = 1;
  ram[3416]  = 1;
  ram[3417]  = 1;
  ram[3418]  = 1;
  ram[3419]  = 1;
  ram[3420]  = 1;
  ram[3421]  = 1;
  ram[3422]  = 1;
  ram[3423]  = 1;
  ram[3424]  = 1;
  ram[3425]  = 1;
  ram[3426]  = 1;
  ram[3427]  = 1;
  ram[3428]  = 1;
  ram[3429]  = 1;
  ram[3430]  = 1;
  ram[3431]  = 1;
  ram[3432]  = 1;
  ram[3433]  = 1;
  ram[3434]  = 1;
  ram[3435]  = 1;
  ram[3436]  = 1;
  ram[3437]  = 1;
  ram[3438]  = 1;
  ram[3439]  = 1;
  ram[3440]  = 1;
  ram[3441]  = 1;
  ram[3442]  = 1;
  ram[3443]  = 1;
  ram[3444]  = 1;
  ram[3445]  = 1;
  ram[3446]  = 1;
  ram[3447]  = 1;
  ram[3448]  = 1;
  ram[3449]  = 1;
  ram[3450]  = 1;
  ram[3451]  = 1;
  ram[3452]  = 1;
  ram[3453]  = 1;
  ram[3454]  = 1;
  ram[3455]  = 1;
  ram[3456]  = 1;
  ram[3457]  = 1;
  ram[3458]  = 1;
  ram[3459]  = 1;
  ram[3460]  = 1;
  ram[3461]  = 1;
  ram[3462]  = 1;
  ram[3463]  = 1;
  ram[3464]  = 1;
  ram[3465]  = 1;
  ram[3466]  = 1;
  ram[3467]  = 1;
  ram[3468]  = 1;
  ram[3469]  = 1;
  ram[3470]  = 1;
  ram[3471]  = 1;
  ram[3472]  = 1;
  ram[3473]  = 1;
  ram[3474]  = 1;
  ram[3475]  = 1;
  ram[3476]  = 1;
  ram[3477]  = 1;
  ram[3478]  = 1;
  ram[3479]  = 1;
  ram[3480]  = 1;
  ram[3481]  = 1;
  ram[3482]  = 1;
  ram[3483]  = 1;
  ram[3484]  = 1;
  ram[3485]  = 1;
  ram[3486]  = 1;
  ram[3487]  = 1;
  ram[3488]  = 1;
  ram[3489]  = 1;
  ram[3490]  = 1;
  ram[3491]  = 1;
  ram[3492]  = 1;
  ram[3493]  = 1;
  ram[3494]  = 1;
  ram[3495]  = 1;
  ram[3496]  = 1;
  ram[3497]  = 1;
  ram[3498]  = 1;
  ram[3499]  = 1;
  ram[3500]  = 1;
  ram[3501]  = 1;
  ram[3502]  = 1;
  ram[3503]  = 1;
  ram[3504]  = 1;
  ram[3505]  = 1;
  ram[3506]  = 1;
  ram[3507]  = 1;
  ram[3508]  = 1;
  ram[3509]  = 1;
  ram[3510]  = 1;
  ram[3511]  = 1;
  ram[3512]  = 1;
  ram[3513]  = 1;
  ram[3514]  = 1;
  ram[3515]  = 1;
  ram[3516]  = 1;
  ram[3517]  = 1;
  ram[3518]  = 1;
  ram[3519]  = 1;
  ram[3520]  = 1;
  ram[3521]  = 1;
  ram[3522]  = 1;
  ram[3523]  = 1;
  ram[3524]  = 1;
  ram[3525]  = 1;
  ram[3526]  = 1;
  ram[3527]  = 1;
  ram[3528]  = 1;
  ram[3529]  = 1;
  ram[3530]  = 1;
  ram[3531]  = 1;
  ram[3532]  = 1;
  ram[3533]  = 1;
  ram[3534]  = 1;
  ram[3535]  = 1;
  ram[3536]  = 1;
  ram[3537]  = 1;
  ram[3538]  = 1;
  ram[3539]  = 1;
  ram[3540]  = 1;
  ram[3541]  = 1;
  ram[3542]  = 1;
  ram[3543]  = 1;
  ram[3544]  = 1;
  ram[3545]  = 1;
  ram[3546]  = 1;
  ram[3547]  = 1;
  ram[3548]  = 1;
  ram[3549]  = 1;
  ram[3550]  = 1;
  ram[3551]  = 1;
  ram[3552]  = 1;
  ram[3553]  = 1;
  ram[3554]  = 1;
  ram[3555]  = 1;
  ram[3556]  = 1;
  ram[3557]  = 1;
  ram[3558]  = 1;
  ram[3559]  = 1;
  ram[3560]  = 1;
  ram[3561]  = 1;
  ram[3562]  = 1;
  ram[3563]  = 1;
  ram[3564]  = 1;
  ram[3565]  = 1;
  ram[3566]  = 1;
  ram[3567]  = 1;
  ram[3568]  = 1;
  ram[3569]  = 1;
  ram[3570]  = 1;
  ram[3571]  = 1;
  ram[3572]  = 1;
  ram[3573]  = 1;
  ram[3574]  = 1;
  ram[3575]  = 1;
  ram[3576]  = 1;
  ram[3577]  = 1;
  ram[3578]  = 1;
  ram[3579]  = 1;
  ram[3580]  = 1;
  ram[3581]  = 1;
  ram[3582]  = 1;
  ram[3583]  = 1;
  ram[3584]  = 1;
  ram[3585]  = 1;
  ram[3586]  = 1;
  ram[3587]  = 1;
  ram[3588]  = 1;
  ram[3589]  = 1;
  ram[3590]  = 1;
  ram[3591]  = 1;
  ram[3592]  = 1;
  ram[3593]  = 1;
  ram[3594]  = 1;
  ram[3595]  = 1;
  ram[3596]  = 1;
  ram[3597]  = 1;
  ram[3598]  = 1;
  ram[3599]  = 1;
  ram[3600]  = 1;
  ram[3601]  = 1;
  ram[3602]  = 1;
  ram[3603]  = 1;
  ram[3604]  = 1;
  ram[3605]  = 1;
  ram[3606]  = 1;
  ram[3607]  = 1;
  ram[3608]  = 1;
  ram[3609]  = 1;
  ram[3610]  = 1;
  ram[3611]  = 1;
  ram[3612]  = 1;
  ram[3613]  = 1;
  ram[3614]  = 1;
  ram[3615]  = 1;
  ram[3616]  = 1;
  ram[3617]  = 1;
  ram[3618]  = 1;
  ram[3619]  = 1;
  ram[3620]  = 1;
  ram[3621]  = 1;
  ram[3622]  = 1;
  ram[3623]  = 1;
  ram[3624]  = 1;
  ram[3625]  = 1;
  ram[3626]  = 1;
  ram[3627]  = 1;
  ram[3628]  = 1;
  ram[3629]  = 1;
  ram[3630]  = 1;
  ram[3631]  = 1;
  ram[3632]  = 1;
  ram[3633]  = 1;
  ram[3634]  = 1;
  ram[3635]  = 1;
  ram[3636]  = 1;
  ram[3637]  = 1;
  ram[3638]  = 1;
  ram[3639]  = 1;
  ram[3640]  = 1;
  ram[3641]  = 1;
  ram[3642]  = 1;
  ram[3643]  = 1;
  ram[3644]  = 1;
  ram[3645]  = 1;
  ram[3646]  = 1;
  ram[3647]  = 1;
  ram[3648]  = 1;
  ram[3649]  = 1;
  ram[3650]  = 1;
  ram[3651]  = 1;
  ram[3652]  = 1;
  ram[3653]  = 1;
  ram[3654]  = 1;
  ram[3655]  = 1;
  ram[3656]  = 1;
  ram[3657]  = 1;
  ram[3658]  = 1;
  ram[3659]  = 1;
  ram[3660]  = 1;
  ram[3661]  = 1;
  ram[3662]  = 1;
  ram[3663]  = 1;
  ram[3664]  = 1;
  ram[3665]  = 1;
  ram[3666]  = 1;
  ram[3667]  = 1;
  ram[3668]  = 1;
  ram[3669]  = 1;
  ram[3670]  = 1;
  ram[3671]  = 1;
  ram[3672]  = 1;
  ram[3673]  = 1;
  ram[3674]  = 1;
  ram[3675]  = 1;
  ram[3676]  = 1;
  ram[3677]  = 1;
  ram[3678]  = 1;
  ram[3679]  = 1;
  ram[3680]  = 1;
  ram[3681]  = 1;
  ram[3682]  = 1;
  ram[3683]  = 1;
  ram[3684]  = 1;
  ram[3685]  = 1;
  ram[3686]  = 1;
  ram[3687]  = 1;
  ram[3688]  = 1;
  ram[3689]  = 1;
  ram[3690]  = 1;
  ram[3691]  = 1;
  ram[3692]  = 1;
  ram[3693]  = 1;
  ram[3694]  = 1;
  ram[3695]  = 1;
  ram[3696]  = 1;
  ram[3697]  = 1;
  ram[3698]  = 1;
  ram[3699]  = 1;
  ram[3700]  = 1;
  ram[3701]  = 1;
  ram[3702]  = 1;
  ram[3703]  = 1;
  ram[3704]  = 1;
  ram[3705]  = 1;
  ram[3706]  = 1;
  ram[3707]  = 1;
  ram[3708]  = 1;
  ram[3709]  = 1;
  ram[3710]  = 1;
  ram[3711]  = 1;
  ram[3712]  = 1;
  ram[3713]  = 1;
  ram[3714]  = 1;
  ram[3715]  = 1;
  ram[3716]  = 1;
  ram[3717]  = 1;
  ram[3718]  = 1;
  ram[3719]  = 1;
  ram[3720]  = 1;
  ram[3721]  = 1;
  ram[3722]  = 1;
  ram[3723]  = 1;
  ram[3724]  = 1;
  ram[3725]  = 1;
  ram[3726]  = 1;
  ram[3727]  = 1;
  ram[3728]  = 1;
  ram[3729]  = 1;
  ram[3730]  = 1;
  ram[3731]  = 1;
  ram[3732]  = 1;
  ram[3733]  = 1;
  ram[3734]  = 1;
  ram[3735]  = 1;
  ram[3736]  = 1;
  ram[3737]  = 1;
  ram[3738]  = 1;
  ram[3739]  = 1;
  ram[3740]  = 1;
  ram[3741]  = 1;
  ram[3742]  = 1;
  ram[3743]  = 1;
  ram[3744]  = 1;
  ram[3745]  = 1;
  ram[3746]  = 1;
  ram[3747]  = 1;
  ram[3748]  = 1;
  ram[3749]  = 1;
  ram[3750]  = 1;
  ram[3751]  = 1;
  ram[3752]  = 1;
  ram[3753]  = 1;
  ram[3754]  = 1;
  ram[3755]  = 1;
  ram[3756]  = 1;
  ram[3757]  = 1;
  ram[3758]  = 1;
  ram[3759]  = 1;
  ram[3760]  = 1;
  ram[3761]  = 1;
  ram[3762]  = 1;
  ram[3763]  = 1;
  ram[3764]  = 1;
  ram[3765]  = 1;
  ram[3766]  = 1;
  ram[3767]  = 1;
  ram[3768]  = 1;
  ram[3769]  = 1;
  ram[3770]  = 1;
  ram[3771]  = 1;
  ram[3772]  = 1;
  ram[3773]  = 1;
  ram[3774]  = 1;
  ram[3775]  = 1;
  ram[3776]  = 1;
  ram[3777]  = 1;
  ram[3778]  = 1;
  ram[3779]  = 1;
  ram[3780]  = 1;
  ram[3781]  = 1;
  ram[3782]  = 1;
  ram[3783]  = 1;
  ram[3784]  = 1;
  ram[3785]  = 1;
  ram[3786]  = 1;
  ram[3787]  = 1;
  ram[3788]  = 1;
  ram[3789]  = 1;
  ram[3790]  = 1;
  ram[3791]  = 1;
  ram[3792]  = 1;
  ram[3793]  = 1;
  ram[3794]  = 1;
  ram[3795]  = 1;
  ram[3796]  = 1;
  ram[3797]  = 1;
  ram[3798]  = 1;
  ram[3799]  = 1;
  ram[3800]  = 1;
  ram[3801]  = 1;
  ram[3802]  = 1;
  ram[3803]  = 1;
  ram[3804]  = 1;
  ram[3805]  = 1;
  ram[3806]  = 1;
  ram[3807]  = 1;
  ram[3808]  = 1;
  ram[3809]  = 1;
  ram[3810]  = 1;
  ram[3811]  = 1;
  ram[3812]  = 1;
  ram[3813]  = 1;
  ram[3814]  = 1;
  ram[3815]  = 1;
  ram[3816]  = 1;
  ram[3817]  = 1;
  ram[3818]  = 1;
  ram[3819]  = 1;
  ram[3820]  = 1;
  ram[3821]  = 1;
  ram[3822]  = 1;
  ram[3823]  = 1;
  ram[3824]  = 1;
  ram[3825]  = 1;
  ram[3826]  = 1;
  ram[3827]  = 1;
  ram[3828]  = 1;
  ram[3829]  = 1;
  ram[3830]  = 1;
  ram[3831]  = 1;
  ram[3832]  = 1;
  ram[3833]  = 1;
  ram[3834]  = 1;
  ram[3835]  = 1;
  ram[3836]  = 1;
  ram[3837]  = 1;
  ram[3838]  = 1;
  ram[3839]  = 1;
  ram[3840]  = 1;
  ram[3841]  = 1;
  ram[3842]  = 1;
  ram[3843]  = 1;
  ram[3844]  = 1;
  ram[3845]  = 1;
  ram[3846]  = 1;
  ram[3847]  = 1;
  ram[3848]  = 1;
  ram[3849]  = 1;
  ram[3850]  = 1;
  ram[3851]  = 1;
  ram[3852]  = 1;
  ram[3853]  = 1;
  ram[3854]  = 1;
  ram[3855]  = 1;
  ram[3856]  = 1;
  ram[3857]  = 1;
  ram[3858]  = 1;
  ram[3859]  = 1;
  ram[3860]  = 1;
  ram[3861]  = 1;
  ram[3862]  = 1;
  ram[3863]  = 1;
  ram[3864]  = 1;
  ram[3865]  = 1;
  ram[3866]  = 1;
  ram[3867]  = 1;
  ram[3868]  = 1;
  ram[3869]  = 1;
  ram[3870]  = 1;
  ram[3871]  = 1;
  ram[3872]  = 1;
  ram[3873]  = 1;
  ram[3874]  = 1;
  ram[3875]  = 1;
  ram[3876]  = 1;
  ram[3877]  = 1;
  ram[3878]  = 1;
  ram[3879]  = 1;
  ram[3880]  = 1;
  ram[3881]  = 1;
  ram[3882]  = 1;
  ram[3883]  = 1;
  ram[3884]  = 1;
  ram[3885]  = 1;
  ram[3886]  = 1;
  ram[3887]  = 1;
  ram[3888]  = 1;
  ram[3889]  = 1;
  ram[3890]  = 1;
  ram[3891]  = 1;
  ram[3892]  = 1;
  ram[3893]  = 1;
  ram[3894]  = 1;
  ram[3895]  = 1;
  ram[3896]  = 1;
  ram[3897]  = 1;
  ram[3898]  = 1;
  ram[3899]  = 1;
  ram[3900]  = 1;
  ram[3901]  = 1;
  ram[3902]  = 1;
  ram[3903]  = 1;
  ram[3904]  = 1;
  ram[3905]  = 1;
  ram[3906]  = 1;
  ram[3907]  = 1;
  ram[3908]  = 1;
  ram[3909]  = 1;
  ram[3910]  = 1;
  ram[3911]  = 1;
  ram[3912]  = 1;
  ram[3913]  = 1;
  ram[3914]  = 1;
  ram[3915]  = 1;
  ram[3916]  = 1;
  ram[3917]  = 1;
  ram[3918]  = 1;
  ram[3919]  = 1;
  ram[3920]  = 1;
  ram[3921]  = 1;
  ram[3922]  = 1;
  ram[3923]  = 1;
  ram[3924]  = 1;
  ram[3925]  = 1;
  ram[3926]  = 1;
  ram[3927]  = 1;
  ram[3928]  = 1;
  ram[3929]  = 1;
  ram[3930]  = 1;
  ram[3931]  = 1;
  ram[3932]  = 1;
  ram[3933]  = 1;
  ram[3934]  = 1;
  ram[3935]  = 1;
  ram[3936]  = 1;
  ram[3937]  = 1;
  ram[3938]  = 1;
  ram[3939]  = 1;
  ram[3940]  = 1;
  ram[3941]  = 1;
  ram[3942]  = 1;
  ram[3943]  = 1;
  ram[3944]  = 1;
  ram[3945]  = 1;
  ram[3946]  = 1;
  ram[3947]  = 1;
  ram[3948]  = 1;
  ram[3949]  = 1;
  ram[3950]  = 1;
  ram[3951]  = 1;
  ram[3952]  = 1;
  ram[3953]  = 1;
  ram[3954]  = 1;
  ram[3955]  = 1;
  ram[3956]  = 1;
  ram[3957]  = 1;
  ram[3958]  = 1;
  ram[3959]  = 1;
  ram[3960]  = 1;
  ram[3961]  = 1;
  ram[3962]  = 1;
  ram[3963]  = 1;
  ram[3964]  = 1;
  ram[3965]  = 1;
  ram[3966]  = 1;
  ram[3967]  = 1;
  ram[3968]  = 1;
  ram[3969]  = 1;
  ram[3970]  = 1;
  ram[3971]  = 1;
  ram[3972]  = 1;
  ram[3973]  = 1;
  ram[3974]  = 1;
  ram[3975]  = 1;
  ram[3976]  = 1;
  ram[3977]  = 1;
  ram[3978]  = 1;
  ram[3979]  = 1;
  ram[3980]  = 1;
  ram[3981]  = 1;
  ram[3982]  = 1;
  ram[3983]  = 1;
  ram[3984]  = 1;
  ram[3985]  = 1;
  ram[3986]  = 1;
  ram[3987]  = 1;
  ram[3988]  = 1;
  ram[3989]  = 1;
  ram[3990]  = 1;
  ram[3991]  = 1;
  ram[3992]  = 1;
  ram[3993]  = 1;
  ram[3994]  = 1;
  ram[3995]  = 1;
  ram[3996]  = 1;
  ram[3997]  = 1;
  ram[3998]  = 1;
  ram[3999]  = 1;
  ram[4000]  = 1;
  ram[4001]  = 1;
  ram[4002]  = 1;
  ram[4003]  = 1;
  ram[4004]  = 1;
  ram[4005]  = 1;
  ram[4006]  = 1;
  ram[4007]  = 1;
  ram[4008]  = 1;
  ram[4009]  = 1;
  ram[4010]  = 1;
  ram[4011]  = 1;
  ram[4012]  = 1;
  ram[4013]  = 1;
  ram[4014]  = 1;
  ram[4015]  = 1;
  ram[4016]  = 1;
  ram[4017]  = 1;
  ram[4018]  = 1;
  ram[4019]  = 1;
  ram[4020]  = 1;
  ram[4021]  = 1;
  ram[4022]  = 1;
  ram[4023]  = 1;
  ram[4024]  = 1;
  ram[4025]  = 1;
  ram[4026]  = 1;
  ram[4027]  = 1;
  ram[4028]  = 1;
  ram[4029]  = 1;
  ram[4030]  = 1;
  ram[4031]  = 1;
  ram[4032]  = 1;
  ram[4033]  = 1;
  ram[4034]  = 1;
  ram[4035]  = 1;
  ram[4036]  = 1;
  ram[4037]  = 1;
  ram[4038]  = 1;
  ram[4039]  = 1;
  ram[4040]  = 1;
  ram[4041]  = 1;
  ram[4042]  = 1;
  ram[4043]  = 1;
  ram[4044]  = 1;
  ram[4045]  = 1;
  ram[4046]  = 1;
  ram[4047]  = 1;
  ram[4048]  = 1;
  ram[4049]  = 1;
  ram[4050]  = 1;
  ram[4051]  = 1;
  ram[4052]  = 1;
  ram[4053]  = 1;
  ram[4054]  = 1;
  ram[4055]  = 1;
  ram[4056]  = 1;
  ram[4057]  = 1;
  ram[4058]  = 1;
  ram[4059]  = 1;
  ram[4060]  = 1;
  ram[4061]  = 1;
  ram[4062]  = 1;
  ram[4063]  = 1;
  ram[4064]  = 1;
  ram[4065]  = 1;
  ram[4066]  = 1;
  ram[4067]  = 1;
  ram[4068]  = 1;
  ram[4069]  = 1;
  ram[4070]  = 1;
  ram[4071]  = 1;
  ram[4072]  = 1;
  ram[4073]  = 1;
  ram[4074]  = 1;
  ram[4075]  = 1;
  ram[4076]  = 1;
  ram[4077]  = 1;
  ram[4078]  = 1;
  ram[4079]  = 1;
  ram[4080]  = 1;
  ram[4081]  = 1;
  ram[4082]  = 1;
  ram[4083]  = 1;
  ram[4084]  = 1;
  ram[4085]  = 1;
  ram[4086]  = 1;
  ram[4087]  = 1;
  ram[4088]  = 1;
  ram[4089]  = 1;
  ram[4090]  = 1;
  ram[4091]  = 1;
  ram[4092]  = 1;
  ram[4093]  = 1;
  ram[4094]  = 1;
  ram[4095]  = 1;
  ram[4096]  = 1;
  ram[4097]  = 1;
  ram[4098]  = 1;
  ram[4099]  = 1;
  ram[4100]  = 1;
  ram[4101]  = 1;
  ram[4102]  = 1;
  ram[4103]  = 1;
  ram[4104]  = 1;
  ram[4105]  = 1;
  ram[4106]  = 1;
  ram[4107]  = 1;
  ram[4108]  = 1;
  ram[4109]  = 1;
  ram[4110]  = 1;
  ram[4111]  = 1;
  ram[4112]  = 1;
  ram[4113]  = 1;
  ram[4114]  = 1;
  ram[4115]  = 1;
  ram[4116]  = 1;
  ram[4117]  = 1;
  ram[4118]  = 1;
  ram[4119]  = 1;
  ram[4120]  = 1;
  ram[4121]  = 1;
  ram[4122]  = 1;
  ram[4123]  = 1;
  ram[4124]  = 1;
  ram[4125]  = 1;
  ram[4126]  = 1;
  ram[4127]  = 1;
  ram[4128]  = 1;
  ram[4129]  = 1;
  ram[4130]  = 1;
  ram[4131]  = 1;
  ram[4132]  = 1;
  ram[4133]  = 1;
  ram[4134]  = 1;
  ram[4135]  = 1;
  ram[4136]  = 1;
  ram[4137]  = 1;
  ram[4138]  = 1;
  ram[4139]  = 1;
  ram[4140]  = 1;
  ram[4141]  = 1;
  ram[4142]  = 1;
  ram[4143]  = 1;
  ram[4144]  = 1;
  ram[4145]  = 1;
  ram[4146]  = 1;
  ram[4147]  = 1;
  ram[4148]  = 1;
  ram[4149]  = 1;
  ram[4150]  = 1;
  ram[4151]  = 1;
  ram[4152]  = 1;
  ram[4153]  = 1;
  ram[4154]  = 1;
  ram[4155]  = 1;
  ram[4156]  = 1;
  ram[4157]  = 1;
  ram[4158]  = 1;
  ram[4159]  = 1;
  ram[4160]  = 1;
  ram[4161]  = 1;
  ram[4162]  = 1;
  ram[4163]  = 1;
  ram[4164]  = 1;
  ram[4165]  = 1;
  ram[4166]  = 1;
  ram[4167]  = 1;
  ram[4168]  = 1;
  ram[4169]  = 1;
  ram[4170]  = 1;
  ram[4171]  = 1;
  ram[4172]  = 1;
  ram[4173]  = 1;
  ram[4174]  = 1;
  ram[4175]  = 1;
  ram[4176]  = 1;
  ram[4177]  = 1;
  ram[4178]  = 1;
  ram[4179]  = 1;
  ram[4180]  = 1;
  ram[4181]  = 1;
  ram[4182]  = 1;
  ram[4183]  = 1;
  ram[4184]  = 1;
  ram[4185]  = 1;
  ram[4186]  = 1;
  ram[4187]  = 1;
  ram[4188]  = 1;
  ram[4189]  = 1;
  ram[4190]  = 1;
  ram[4191]  = 1;
  ram[4192]  = 1;
  ram[4193]  = 1;
  ram[4194]  = 1;
  ram[4195]  = 1;
  ram[4196]  = 1;
  ram[4197]  = 1;
  ram[4198]  = 1;
  ram[4199]  = 1;
  ram[4200]  = 1;
  ram[4201]  = 1;
  ram[4202]  = 1;
  ram[4203]  = 1;
  ram[4204]  = 1;
  ram[4205]  = 1;
  ram[4206]  = 1;
  ram[4207]  = 1;
  ram[4208]  = 1;
  ram[4209]  = 1;
  ram[4210]  = 1;
  ram[4211]  = 1;
  ram[4212]  = 1;
  ram[4213]  = 1;
  ram[4214]  = 1;
  ram[4215]  = 1;
  ram[4216]  = 1;
  ram[4217]  = 1;
  ram[4218]  = 1;
  ram[4219]  = 1;
  ram[4220]  = 1;
  ram[4221]  = 1;
  ram[4222]  = 1;
  ram[4223]  = 1;
  ram[4224]  = 1;
  ram[4225]  = 1;
  ram[4226]  = 1;
  ram[4227]  = 1;
  ram[4228]  = 1;
  ram[4229]  = 1;
  ram[4230]  = 1;
  ram[4231]  = 1;
  ram[4232]  = 1;
  ram[4233]  = 1;
  ram[4234]  = 1;
  ram[4235]  = 1;
  ram[4236]  = 1;
  ram[4237]  = 1;
  ram[4238]  = 1;
  ram[4239]  = 1;
  ram[4240]  = 1;
  ram[4241]  = 1;
  ram[4242]  = 1;
  ram[4243]  = 1;
  ram[4244]  = 1;
  ram[4245]  = 1;
  ram[4246]  = 1;
  ram[4247]  = 1;
  ram[4248]  = 1;
  ram[4249]  = 1;
  ram[4250]  = 1;
  ram[4251]  = 1;
  ram[4252]  = 1;
  ram[4253]  = 1;
  ram[4254]  = 1;
  ram[4255]  = 1;
  ram[4256]  = 1;
  ram[4257]  = 1;
  ram[4258]  = 1;
  ram[4259]  = 1;
  ram[4260]  = 1;
  ram[4261]  = 1;
  ram[4262]  = 1;
  ram[4263]  = 1;
  ram[4264]  = 1;
  ram[4265]  = 1;
  ram[4266]  = 1;
  ram[4267]  = 1;
  ram[4268]  = 1;
  ram[4269]  = 1;
  ram[4270]  = 1;
  ram[4271]  = 1;
  ram[4272]  = 1;
  ram[4273]  = 1;
  ram[4274]  = 1;
  ram[4275]  = 1;
  ram[4276]  = 1;
  ram[4277]  = 1;
  ram[4278]  = 1;
  ram[4279]  = 1;
  ram[4280]  = 1;
  ram[4281]  = 1;
  ram[4282]  = 1;
  ram[4283]  = 1;
  ram[4284]  = 1;
  ram[4285]  = 1;
  ram[4286]  = 1;
  ram[4287]  = 1;
  ram[4288]  = 1;
  ram[4289]  = 1;
  ram[4290]  = 1;
  ram[4291]  = 1;
  ram[4292]  = 1;
  ram[4293]  = 1;
  ram[4294]  = 1;
  ram[4295]  = 1;
  ram[4296]  = 1;
  ram[4297]  = 1;
  ram[4298]  = 1;
  ram[4299]  = 1;
  ram[4300]  = 1;
  ram[4301]  = 1;
  ram[4302]  = 1;
  ram[4303]  = 1;
  ram[4304]  = 1;
  ram[4305]  = 1;
  ram[4306]  = 1;
  ram[4307]  = 1;
  ram[4308]  = 1;
  ram[4309]  = 1;
  ram[4310]  = 1;
  ram[4311]  = 1;
  ram[4312]  = 1;
  ram[4313]  = 1;
  ram[4314]  = 1;
  ram[4315]  = 1;
  ram[4316]  = 1;
  ram[4317]  = 1;
  ram[4318]  = 1;
  ram[4319]  = 1;
  ram[4320]  = 1;
  ram[4321]  = 1;
  ram[4322]  = 1;
  ram[4323]  = 1;
  ram[4324]  = 1;
  ram[4325]  = 1;
  ram[4326]  = 1;
  ram[4327]  = 1;
  ram[4328]  = 1;
  ram[4329]  = 1;
  ram[4330]  = 1;
  ram[4331]  = 1;
  ram[4332]  = 1;
  ram[4333]  = 1;
  ram[4334]  = 1;
  ram[4335]  = 1;
  ram[4336]  = 1;
  ram[4337]  = 1;
  ram[4338]  = 1;
  ram[4339]  = 1;
  ram[4340]  = 1;
  ram[4341]  = 1;
  ram[4342]  = 1;
  ram[4343]  = 1;
  ram[4344]  = 1;
  ram[4345]  = 1;
  ram[4346]  = 1;
  ram[4347]  = 1;
  ram[4348]  = 1;
  ram[4349]  = 1;
  ram[4350]  = 1;
  ram[4351]  = 1;
  ram[4352]  = 1;
  ram[4353]  = 1;
  ram[4354]  = 1;
  ram[4355]  = 1;
  ram[4356]  = 1;
  ram[4357]  = 1;
  ram[4358]  = 1;
  ram[4359]  = 1;
  ram[4360]  = 1;
  ram[4361]  = 1;
  ram[4362]  = 1;
  ram[4363]  = 1;
  ram[4364]  = 1;
  ram[4365]  = 1;
  ram[4366]  = 1;
  ram[4367]  = 1;
  ram[4368]  = 1;
  ram[4369]  = 1;
  ram[4370]  = 1;
  ram[4371]  = 1;
  ram[4372]  = 1;
  ram[4373]  = 1;
  ram[4374]  = 1;
  ram[4375]  = 1;
  ram[4376]  = 1;
  ram[4377]  = 1;
  ram[4378]  = 1;
  ram[4379]  = 1;
  ram[4380]  = 1;
  ram[4381]  = 1;
  ram[4382]  = 1;
  ram[4383]  = 1;
  ram[4384]  = 1;
  ram[4385]  = 1;
  ram[4386]  = 1;
  ram[4387]  = 1;
  ram[4388]  = 1;
  ram[4389]  = 1;
  ram[4390]  = 1;
  ram[4391]  = 1;
  ram[4392]  = 1;
  ram[4393]  = 1;
  ram[4394]  = 1;
  ram[4395]  = 1;
  ram[4396]  = 1;
  ram[4397]  = 1;
  ram[4398]  = 1;
  ram[4399]  = 1;
  ram[4400]  = 1;
  ram[4401]  = 1;
  ram[4402]  = 1;
  ram[4403]  = 1;
  ram[4404]  = 1;
  ram[4405]  = 1;
  ram[4406]  = 1;
  ram[4407]  = 1;
  ram[4408]  = 1;
  ram[4409]  = 1;
  ram[4410]  = 1;
  ram[4411]  = 1;
  ram[4412]  = 1;
  ram[4413]  = 1;
  ram[4414]  = 1;
  ram[4415]  = 1;
  ram[4416]  = 1;
  ram[4417]  = 1;
  ram[4418]  = 1;
  ram[4419]  = 1;
  ram[4420]  = 1;
  ram[4421]  = 1;
  ram[4422]  = 1;
  ram[4423]  = 1;
  ram[4424]  = 1;
  ram[4425]  = 1;
  ram[4426]  = 1;
  ram[4427]  = 1;
  ram[4428]  = 1;
  ram[4429]  = 1;
  ram[4430]  = 1;
  ram[4431]  = 1;
  ram[4432]  = 1;
  ram[4433]  = 1;
  ram[4434]  = 1;
  ram[4435]  = 1;
  ram[4436]  = 1;
  ram[4437]  = 1;
  ram[4438]  = 1;
  ram[4439]  = 1;
  ram[4440]  = 1;
  ram[4441]  = 1;
  ram[4442]  = 1;
  ram[4443]  = 1;
  ram[4444]  = 1;
  ram[4445]  = 1;
  ram[4446]  = 1;
  ram[4447]  = 1;
  ram[4448]  = 1;
  ram[4449]  = 1;
  ram[4450]  = 1;
  ram[4451]  = 1;
  ram[4452]  = 1;
  ram[4453]  = 1;
  ram[4454]  = 1;
  ram[4455]  = 1;
  ram[4456]  = 1;
  ram[4457]  = 1;
  ram[4458]  = 1;
  ram[4459]  = 1;
  ram[4460]  = 1;
  ram[4461]  = 1;
  ram[4462]  = 1;
  ram[4463]  = 1;
  ram[4464]  = 1;
  ram[4465]  = 1;
  ram[4466]  = 1;
  ram[4467]  = 1;
  ram[4468]  = 1;
  ram[4469]  = 1;
  ram[4470]  = 1;
  ram[4471]  = 1;
  ram[4472]  = 1;
  ram[4473]  = 1;
  ram[4474]  = 1;
  ram[4475]  = 1;
  ram[4476]  = 1;
  ram[4477]  = 1;
  ram[4478]  = 1;
  ram[4479]  = 1;
  ram[4480]  = 1;
  ram[4481]  = 1;
  ram[4482]  = 1;
  ram[4483]  = 1;
  ram[4484]  = 1;
  ram[4485]  = 1;
  ram[4486]  = 1;
  ram[4487]  = 1;
  ram[4488]  = 1;
  ram[4489]  = 1;
  ram[4490]  = 1;
  ram[4491]  = 1;
  ram[4492]  = 1;
  ram[4493]  = 1;
  ram[4494]  = 1;
  ram[4495]  = 1;
  ram[4496]  = 1;
  ram[4497]  = 1;
  ram[4498]  = 1;
  ram[4499]  = 1;
  ram[4500]  = 1;
  ram[4501]  = 1;
  ram[4502]  = 1;
  ram[4503]  = 1;
  ram[4504]  = 1;
  ram[4505]  = 1;
  ram[4506]  = 1;
  ram[4507]  = 1;
  ram[4508]  = 1;
  ram[4509]  = 1;
  ram[4510]  = 1;
  ram[4511]  = 1;
  ram[4512]  = 1;
  ram[4513]  = 1;
  ram[4514]  = 1;
  ram[4515]  = 1;
  ram[4516]  = 1;
  ram[4517]  = 1;
  ram[4518]  = 1;
  ram[4519]  = 1;
  ram[4520]  = 1;
  ram[4521]  = 1;
  ram[4522]  = 1;
  ram[4523]  = 1;
  ram[4524]  = 1;
  ram[4525]  = 1;
  ram[4526]  = 1;
  ram[4527]  = 1;
  ram[4528]  = 1;
  ram[4529]  = 1;
  ram[4530]  = 1;
  ram[4531]  = 1;
  ram[4532]  = 1;
  ram[4533]  = 1;
  ram[4534]  = 1;
  ram[4535]  = 1;
  ram[4536]  = 1;
  ram[4537]  = 1;
  ram[4538]  = 1;
  ram[4539]  = 1;
  ram[4540]  = 1;
  ram[4541]  = 1;
  ram[4542]  = 1;
  ram[4543]  = 1;
  ram[4544]  = 1;
  ram[4545]  = 1;
  ram[4546]  = 1;
  ram[4547]  = 1;
  ram[4548]  = 1;
  ram[4549]  = 1;
  ram[4550]  = 1;
  ram[4551]  = 1;
  ram[4552]  = 1;
  ram[4553]  = 1;
  ram[4554]  = 1;
  ram[4555]  = 1;
  ram[4556]  = 1;
  ram[4557]  = 1;
  ram[4558]  = 1;
  ram[4559]  = 1;
  ram[4560]  = 1;
  ram[4561]  = 1;
  ram[4562]  = 1;
  ram[4563]  = 1;
  ram[4564]  = 1;
  ram[4565]  = 1;
  ram[4566]  = 1;
  ram[4567]  = 1;
  ram[4568]  = 1;
  ram[4569]  = 1;
  ram[4570]  = 1;
  ram[4571]  = 1;
  ram[4572]  = 1;
  ram[4573]  = 1;
  ram[4574]  = 1;
  ram[4575]  = 1;
  ram[4576]  = 1;
  ram[4577]  = 1;
  ram[4578]  = 1;
  ram[4579]  = 1;
  ram[4580]  = 1;
  ram[4581]  = 1;
  ram[4582]  = 1;
  ram[4583]  = 1;
  ram[4584]  = 1;
  ram[4585]  = 1;
  ram[4586]  = 1;
  ram[4587]  = 1;
  ram[4588]  = 1;
  ram[4589]  = 1;
  ram[4590]  = 1;
  ram[4591]  = 1;
  ram[4592]  = 1;
  ram[4593]  = 1;
  ram[4594]  = 1;
  ram[4595]  = 1;
  ram[4596]  = 1;
  ram[4597]  = 1;
  ram[4598]  = 1;
  ram[4599]  = 1;
  ram[4600]  = 1;
  ram[4601]  = 1;
  ram[4602]  = 1;
  ram[4603]  = 1;
  ram[4604]  = 1;
  ram[4605]  = 1;
  ram[4606]  = 1;
  ram[4607]  = 1;
  ram[4608]  = 1;
  ram[4609]  = 1;
  ram[4610]  = 1;
  ram[4611]  = 1;
  ram[4612]  = 1;
  ram[4613]  = 1;
  ram[4614]  = 1;
  ram[4615]  = 1;
  ram[4616]  = 1;
  ram[4617]  = 1;
  ram[4618]  = 1;
  ram[4619]  = 1;
  ram[4620]  = 1;
  ram[4621]  = 1;
  ram[4622]  = 1;
  ram[4623]  = 1;
  ram[4624]  = 1;
  ram[4625]  = 1;
  ram[4626]  = 1;
  ram[4627]  = 1;
  ram[4628]  = 1;
  ram[4629]  = 1;
  ram[4630]  = 1;
  ram[4631]  = 1;
  ram[4632]  = 1;
  ram[4633]  = 1;
  ram[4634]  = 1;
  ram[4635]  = 1;
  ram[4636]  = 1;
  ram[4637]  = 1;
  ram[4638]  = 1;
  ram[4639]  = 1;
  ram[4640]  = 1;
  ram[4641]  = 1;
  ram[4642]  = 1;
  ram[4643]  = 1;
  ram[4644]  = 1;
  ram[4645]  = 1;
  ram[4646]  = 1;
  ram[4647]  = 1;
  ram[4648]  = 1;
  ram[4649]  = 1;
  ram[4650]  = 1;
  ram[4651]  = 1;
  ram[4652]  = 1;
  ram[4653]  = 1;
  ram[4654]  = 1;
  ram[4655]  = 1;
  ram[4656]  = 1;
  ram[4657]  = 1;
  ram[4658]  = 1;
  ram[4659]  = 1;
  ram[4660]  = 1;
  ram[4661]  = 1;
  ram[4662]  = 1;
  ram[4663]  = 1;
  ram[4664]  = 1;
  ram[4665]  = 1;
  ram[4666]  = 1;
  ram[4667]  = 1;
  ram[4668]  = 1;
  ram[4669]  = 1;
  ram[4670]  = 1;
  ram[4671]  = 1;
  ram[4672]  = 1;
  ram[4673]  = 1;
  ram[4674]  = 1;
  ram[4675]  = 1;
  ram[4676]  = 1;
  ram[4677]  = 1;
  ram[4678]  = 1;
  ram[4679]  = 1;
  ram[4680]  = 1;
  ram[4681]  = 1;
  ram[4682]  = 1;
  ram[4683]  = 1;
  ram[4684]  = 1;
  ram[4685]  = 1;
  ram[4686]  = 1;
  ram[4687]  = 1;
  ram[4688]  = 1;
  ram[4689]  = 1;
  ram[4690]  = 1;
  ram[4691]  = 1;
  ram[4692]  = 1;
  ram[4693]  = 1;
  ram[4694]  = 1;
  ram[4695]  = 1;
  ram[4696]  = 1;
  ram[4697]  = 1;
  ram[4698]  = 1;
  ram[4699]  = 1;
  ram[4700]  = 1;
  ram[4701]  = 1;
  ram[4702]  = 1;
  ram[4703]  = 1;
  ram[4704]  = 1;
  ram[4705]  = 1;
  ram[4706]  = 1;
  ram[4707]  = 1;
  ram[4708]  = 1;
  ram[4709]  = 1;
  ram[4710]  = 1;
  ram[4711]  = 1;
  ram[4712]  = 1;
  ram[4713]  = 1;
  ram[4714]  = 1;
  ram[4715]  = 1;
  ram[4716]  = 1;
  ram[4717]  = 1;
  ram[4718]  = 1;
  ram[4719]  = 1;
  ram[4720]  = 1;
  ram[4721]  = 1;
  ram[4722]  = 1;
  ram[4723]  = 1;
  ram[4724]  = 1;
  ram[4725]  = 1;
  ram[4726]  = 1;
  ram[4727]  = 1;
  ram[4728]  = 1;
  ram[4729]  = 1;
  ram[4730]  = 1;
  ram[4731]  = 1;
  ram[4732]  = 1;
  ram[4733]  = 1;
  ram[4734]  = 1;
  ram[4735]  = 1;
  ram[4736]  = 1;
  ram[4737]  = 1;
  ram[4738]  = 1;
  ram[4739]  = 1;
  ram[4740]  = 1;
  ram[4741]  = 1;
  ram[4742]  = 1;
  ram[4743]  = 1;
  ram[4744]  = 1;
  ram[4745]  = 1;
  ram[4746]  = 1;
  ram[4747]  = 1;
  ram[4748]  = 1;
  ram[4749]  = 1;
  ram[4750]  = 1;
  ram[4751]  = 1;
  ram[4752]  = 1;
  ram[4753]  = 1;
  ram[4754]  = 1;
  ram[4755]  = 1;
  ram[4756]  = 1;
  ram[4757]  = 1;
  ram[4758]  = 1;
  ram[4759]  = 1;
  ram[4760]  = 1;
  ram[4761]  = 1;
  ram[4762]  = 1;
  ram[4763]  = 1;
  ram[4764]  = 1;
  ram[4765]  = 1;
  ram[4766]  = 1;
  ram[4767]  = 1;
  ram[4768]  = 1;
  ram[4769]  = 1;
  ram[4770]  = 1;
  ram[4771]  = 1;
  ram[4772]  = 1;
  ram[4773]  = 1;
  ram[4774]  = 1;
  ram[4775]  = 1;
  ram[4776]  = 1;
  ram[4777]  = 1;
  ram[4778]  = 1;
  ram[4779]  = 1;
  ram[4780]  = 1;
  ram[4781]  = 1;
  ram[4782]  = 1;
  ram[4783]  = 1;
  ram[4784]  = 1;
  ram[4785]  = 1;
  ram[4786]  = 1;
  ram[4787]  = 1;
  ram[4788]  = 1;
  ram[4789]  = 1;
  ram[4790]  = 1;
  ram[4791]  = 1;
  ram[4792]  = 1;
  ram[4793]  = 1;
  ram[4794]  = 1;
  ram[4795]  = 1;
  ram[4796]  = 1;
  ram[4797]  = 1;
  ram[4798]  = 1;
  ram[4799]  = 1;
  ram[4800]  = 1;
  ram[4801]  = 1;
  ram[4802]  = 1;
  ram[4803]  = 1;
  ram[4804]  = 1;
  ram[4805]  = 1;
  ram[4806]  = 1;
  ram[4807]  = 1;
  ram[4808]  = 1;
  ram[4809]  = 1;
  ram[4810]  = 1;
  ram[4811]  = 1;
  ram[4812]  = 1;
  ram[4813]  = 1;
  ram[4814]  = 1;
  ram[4815]  = 1;
  ram[4816]  = 1;
  ram[4817]  = 1;
  ram[4818]  = 1;
  ram[4819]  = 1;
  ram[4820]  = 1;
  ram[4821]  = 1;
  ram[4822]  = 1;
  ram[4823]  = 1;
  ram[4824]  = 1;
  ram[4825]  = 1;
  ram[4826]  = 1;
  ram[4827]  = 1;
  ram[4828]  = 1;
  ram[4829]  = 1;
  ram[4830]  = 1;
  ram[4831]  = 1;
  ram[4832]  = 1;
  ram[4833]  = 1;
  ram[4834]  = 1;
  ram[4835]  = 1;
  ram[4836]  = 1;
  ram[4837]  = 1;
  ram[4838]  = 1;
  ram[4839]  = 1;
  ram[4840]  = 1;
  ram[4841]  = 1;
  ram[4842]  = 1;
  ram[4843]  = 1;
  ram[4844]  = 1;
  ram[4845]  = 1;
  ram[4846]  = 1;
  ram[4847]  = 1;
  ram[4848]  = 1;
  ram[4849]  = 1;
  ram[4850]  = 1;
  ram[4851]  = 1;
  ram[4852]  = 1;
  ram[4853]  = 1;
  ram[4854]  = 1;
  ram[4855]  = 1;
  ram[4856]  = 1;
  ram[4857]  = 1;
  ram[4858]  = 1;
  ram[4859]  = 1;
  ram[4860]  = 1;
  ram[4861]  = 1;
  ram[4862]  = 1;
  ram[4863]  = 1;
  ram[4864]  = 1;
  ram[4865]  = 1;
  ram[4866]  = 1;
  ram[4867]  = 1;
  ram[4868]  = 1;
  ram[4869]  = 1;
  ram[4870]  = 1;
  ram[4871]  = 1;
  ram[4872]  = 1;
  ram[4873]  = 1;
  ram[4874]  = 1;
  ram[4875]  = 1;
  ram[4876]  = 1;
  ram[4877]  = 1;
  ram[4878]  = 1;
  ram[4879]  = 1;
  ram[4880]  = 1;
  ram[4881]  = 1;
  ram[4882]  = 1;
  ram[4883]  = 1;
  ram[4884]  = 1;
  ram[4885]  = 1;
  ram[4886]  = 1;
  ram[4887]  = 1;
  ram[4888]  = 1;
  ram[4889]  = 1;
  ram[4890]  = 1;
  ram[4891]  = 1;
  ram[4892]  = 1;
  ram[4893]  = 1;
  ram[4894]  = 1;
  ram[4895]  = 1;
  ram[4896]  = 1;
  ram[4897]  = 1;
  ram[4898]  = 1;
  ram[4899]  = 1;
  ram[4900]  = 1;
  ram[4901]  = 1;
  ram[4902]  = 1;
  ram[4903]  = 1;
  ram[4904]  = 1;
  ram[4905]  = 1;
  ram[4906]  = 1;
  ram[4907]  = 1;
  ram[4908]  = 1;
  ram[4909]  = 1;
  ram[4910]  = 1;
  ram[4911]  = 1;
  ram[4912]  = 1;
  ram[4913]  = 1;
  ram[4914]  = 1;
  ram[4915]  = 1;
  ram[4916]  = 1;
  ram[4917]  = 1;
  ram[4918]  = 1;
  ram[4919]  = 1;
  ram[4920]  = 1;
  ram[4921]  = 1;
  ram[4922]  = 1;
  ram[4923]  = 1;
  ram[4924]  = 1;
  ram[4925]  = 1;
  ram[4926]  = 1;
  ram[4927]  = 1;
  ram[4928]  = 1;
  ram[4929]  = 1;
  ram[4930]  = 1;
  ram[4931]  = 1;
  ram[4932]  = 1;
  ram[4933]  = 1;
  ram[4934]  = 1;
  ram[4935]  = 1;
  ram[4936]  = 1;
  ram[4937]  = 1;
  ram[4938]  = 1;
  ram[4939]  = 1;
  ram[4940]  = 1;
  ram[4941]  = 1;
  ram[4942]  = 1;
  ram[4943]  = 1;
  ram[4944]  = 1;
  ram[4945]  = 1;
  ram[4946]  = 1;
  ram[4947]  = 1;
  ram[4948]  = 1;
  ram[4949]  = 1;
  ram[4950]  = 1;
  ram[4951]  = 1;
  ram[4952]  = 1;
  ram[4953]  = 1;
  ram[4954]  = 1;
  ram[4955]  = 1;
  ram[4956]  = 1;
  ram[4957]  = 1;
  ram[4958]  = 1;
  ram[4959]  = 1;
  ram[4960]  = 1;
  ram[4961]  = 1;
  ram[4962]  = 1;
  ram[4963]  = 1;
  ram[4964]  = 1;
  ram[4965]  = 1;
  ram[4966]  = 1;
  ram[4967]  = 1;
  ram[4968]  = 1;
  ram[4969]  = 1;
  ram[4970]  = 1;
  ram[4971]  = 1;
  ram[4972]  = 1;
  ram[4973]  = 1;
  ram[4974]  = 1;
  ram[4975]  = 1;
  ram[4976]  = 1;
  ram[4977]  = 1;
  ram[4978]  = 1;
  ram[4979]  = 1;
  ram[4980]  = 1;
  ram[4981]  = 1;
  ram[4982]  = 1;
  ram[4983]  = 1;
  ram[4984]  = 1;
  ram[4985]  = 1;
  ram[4986]  = 1;
  ram[4987]  = 1;
  ram[4988]  = 1;
  ram[4989]  = 1;
  ram[4990]  = 1;
  ram[4991]  = 1;
  ram[4992]  = 1;
  ram[4993]  = 1;
  ram[4994]  = 1;
  ram[4995]  = 1;
  ram[4996]  = 1;
  ram[4997]  = 1;
  ram[4998]  = 1;
  ram[4999]  = 1;
  ram[5000]  = 1;
  ram[5001]  = 1;
  ram[5002]  = 1;
  ram[5003]  = 1;
  ram[5004]  = 1;
  ram[5005]  = 1;
  ram[5006]  = 1;
  ram[5007]  = 1;
  ram[5008]  = 1;
  ram[5009]  = 1;
  ram[5010]  = 1;
  ram[5011]  = 1;
  ram[5012]  = 1;
  ram[5013]  = 1;
  ram[5014]  = 1;
  ram[5015]  = 1;
  ram[5016]  = 1;
  ram[5017]  = 1;
  ram[5018]  = 1;
  ram[5019]  = 1;
  ram[5020]  = 1;
  ram[5021]  = 1;
  ram[5022]  = 1;
  ram[5023]  = 1;
  ram[5024]  = 1;
  ram[5025]  = 1;
  ram[5026]  = 1;
  ram[5027]  = 1;
  ram[5028]  = 1;
  ram[5029]  = 1;
  ram[5030]  = 1;
  ram[5031]  = 1;
  ram[5032]  = 1;
  ram[5033]  = 1;
  ram[5034]  = 1;
  ram[5035]  = 1;
  ram[5036]  = 1;
  ram[5037]  = 1;
  ram[5038]  = 1;
  ram[5039]  = 1;
  ram[5040]  = 1;
  ram[5041]  = 1;
  ram[5042]  = 1;
  ram[5043]  = 1;
  ram[5044]  = 1;
  ram[5045]  = 1;
  ram[5046]  = 1;
  ram[5047]  = 1;
  ram[5048]  = 1;
  ram[5049]  = 1;
  ram[5050]  = 1;
  ram[5051]  = 1;
  ram[5052]  = 1;
  ram[5053]  = 1;
  ram[5054]  = 1;
  ram[5055]  = 1;
  ram[5056]  = 1;
  ram[5057]  = 1;
  ram[5058]  = 1;
  ram[5059]  = 1;
  ram[5060]  = 1;
  ram[5061]  = 1;
  ram[5062]  = 1;
  ram[5063]  = 1;
  ram[5064]  = 1;
  ram[5065]  = 1;
  ram[5066]  = 1;
  ram[5067]  = 1;
  ram[5068]  = 1;
  ram[5069]  = 1;
  ram[5070]  = 1;
  ram[5071]  = 1;
  ram[5072]  = 1;
  ram[5073]  = 1;
  ram[5074]  = 1;
  ram[5075]  = 1;
  ram[5076]  = 1;
  ram[5077]  = 1;
  ram[5078]  = 1;
  ram[5079]  = 1;
  ram[5080]  = 1;
  ram[5081]  = 1;
  ram[5082]  = 1;
  ram[5083]  = 1;
  ram[5084]  = 1;
  ram[5085]  = 1;
  ram[5086]  = 1;
  ram[5087]  = 1;
  ram[5088]  = 1;
  ram[5089]  = 1;
  ram[5090]  = 1;
  ram[5091]  = 1;
  ram[5092]  = 1;
  ram[5093]  = 1;
  ram[5094]  = 1;
  ram[5095]  = 1;
  ram[5096]  = 1;
  ram[5097]  = 1;
  ram[5098]  = 1;
  ram[5099]  = 1;
  ram[5100]  = 1;
  ram[5101]  = 1;
  ram[5102]  = 1;
  ram[5103]  = 1;
  ram[5104]  = 1;
  ram[5105]  = 1;
  ram[5106]  = 1;
  ram[5107]  = 1;
  ram[5108]  = 1;
  ram[5109]  = 1;
  ram[5110]  = 1;
  ram[5111]  = 1;
  ram[5112]  = 1;
  ram[5113]  = 1;
  ram[5114]  = 1;
  ram[5115]  = 1;
  ram[5116]  = 1;
  ram[5117]  = 1;
  ram[5118]  = 1;
  ram[5119]  = 1;
  ram[5120]  = 1;
  ram[5121]  = 1;
  ram[5122]  = 1;
  ram[5123]  = 1;
  ram[5124]  = 1;
  ram[5125]  = 1;
  ram[5126]  = 1;
  ram[5127]  = 1;
  ram[5128]  = 1;
  ram[5129]  = 1;
  ram[5130]  = 1;
  ram[5131]  = 1;
  ram[5132]  = 1;
  ram[5133]  = 1;
  ram[5134]  = 1;
  ram[5135]  = 1;
  ram[5136]  = 1;
  ram[5137]  = 1;
  ram[5138]  = 1;
  ram[5139]  = 1;
  ram[5140]  = 1;
  ram[5141]  = 1;
  ram[5142]  = 1;
  ram[5143]  = 1;
  ram[5144]  = 1;
  ram[5145]  = 1;
  ram[5146]  = 1;
  ram[5147]  = 1;
  ram[5148]  = 1;
  ram[5149]  = 1;
  ram[5150]  = 1;
  ram[5151]  = 1;
  ram[5152]  = 1;
  ram[5153]  = 1;
  ram[5154]  = 1;
  ram[5155]  = 1;
  ram[5156]  = 1;
  ram[5157]  = 1;
  ram[5158]  = 1;
  ram[5159]  = 1;
  ram[5160]  = 1;
  ram[5161]  = 1;
  ram[5162]  = 1;
  ram[5163]  = 1;
  ram[5164]  = 1;
  ram[5165]  = 1;
  ram[5166]  = 1;
  ram[5167]  = 1;
  ram[5168]  = 1;
  ram[5169]  = 1;
  ram[5170]  = 1;
  ram[5171]  = 1;
  ram[5172]  = 1;
  ram[5173]  = 1;
  ram[5174]  = 1;
  ram[5175]  = 1;
  ram[5176]  = 1;
  ram[5177]  = 1;
  ram[5178]  = 1;
  ram[5179]  = 1;
  ram[5180]  = 1;
  ram[5181]  = 1;
  ram[5182]  = 1;
  ram[5183]  = 1;
  ram[5184]  = 1;
  ram[5185]  = 1;
  ram[5186]  = 1;
  ram[5187]  = 1;
  ram[5188]  = 1;
  ram[5189]  = 1;
  ram[5190]  = 1;
  ram[5191]  = 1;
  ram[5192]  = 1;
  ram[5193]  = 1;
  ram[5194]  = 1;
  ram[5195]  = 1;
  ram[5196]  = 1;
  ram[5197]  = 1;
  ram[5198]  = 1;
  ram[5199]  = 1;
  ram[5200]  = 1;
  ram[5201]  = 1;
  ram[5202]  = 1;
  ram[5203]  = 1;
  ram[5204]  = 1;
  ram[5205]  = 1;
  ram[5206]  = 1;
  ram[5207]  = 1;
  ram[5208]  = 1;
  ram[5209]  = 1;
  ram[5210]  = 1;
  ram[5211]  = 1;
  ram[5212]  = 1;
  ram[5213]  = 1;
  ram[5214]  = 1;
  ram[5215]  = 1;
  ram[5216]  = 1;
  ram[5217]  = 1;
  ram[5218]  = 1;
  ram[5219]  = 1;
  ram[5220]  = 1;
  ram[5221]  = 1;
  ram[5222]  = 1;
  ram[5223]  = 1;
  ram[5224]  = 1;
  ram[5225]  = 1;
  ram[5226]  = 1;
  ram[5227]  = 1;
  ram[5228]  = 1;
  ram[5229]  = 1;
  ram[5230]  = 1;
  ram[5231]  = 1;
  ram[5232]  = 1;
  ram[5233]  = 1;
  ram[5234]  = 1;
  ram[5235]  = 1;
  ram[5236]  = 1;
  ram[5237]  = 1;
  ram[5238]  = 1;
  ram[5239]  = 1;
  ram[5240]  = 1;
  ram[5241]  = 1;
  ram[5242]  = 1;
  ram[5243]  = 1;
  ram[5244]  = 1;
  ram[5245]  = 1;
  ram[5246]  = 1;
  ram[5247]  = 1;
  ram[5248]  = 1;
  ram[5249]  = 1;
  ram[5250]  = 1;
  ram[5251]  = 1;
  ram[5252]  = 1;
  ram[5253]  = 1;
  ram[5254]  = 1;
  ram[5255]  = 1;
  ram[5256]  = 1;
  ram[5257]  = 1;
  ram[5258]  = 1;
  ram[5259]  = 1;
  ram[5260]  = 1;
  ram[5261]  = 1;
  ram[5262]  = 1;
  ram[5263]  = 1;
  ram[5264]  = 1;
  ram[5265]  = 1;
  ram[5266]  = 1;
  ram[5267]  = 1;
  ram[5268]  = 1;
  ram[5269]  = 1;
  ram[5270]  = 1;
  ram[5271]  = 1;
  ram[5272]  = 1;
  ram[5273]  = 1;
  ram[5274]  = 1;
  ram[5275]  = 1;
  ram[5276]  = 1;
  ram[5277]  = 1;
  ram[5278]  = 1;
  ram[5279]  = 1;
  ram[5280]  = 1;
  ram[5281]  = 1;
  ram[5282]  = 1;
  ram[5283]  = 1;
  ram[5284]  = 1;
  ram[5285]  = 1;
  ram[5286]  = 1;
  ram[5287]  = 1;
  ram[5288]  = 1;
  ram[5289]  = 1;
  ram[5290]  = 1;
  ram[5291]  = 1;
  ram[5292]  = 1;
  ram[5293]  = 1;
  ram[5294]  = 1;
  ram[5295]  = 1;
  ram[5296]  = 1;
  ram[5297]  = 1;
  ram[5298]  = 1;
  ram[5299]  = 1;
  ram[5300]  = 1;
  ram[5301]  = 1;
  ram[5302]  = 1;
  ram[5303]  = 1;
  ram[5304]  = 1;
  ram[5305]  = 1;
  ram[5306]  = 1;
  ram[5307]  = 1;
  ram[5308]  = 1;
  ram[5309]  = 1;
  ram[5310]  = 1;
  ram[5311]  = 1;
  ram[5312]  = 1;
  ram[5313]  = 1;
  ram[5314]  = 1;
  ram[5315]  = 1;
  ram[5316]  = 1;
  ram[5317]  = 1;
  ram[5318]  = 1;
  ram[5319]  = 1;
  ram[5320]  = 1;
  ram[5321]  = 1;
  ram[5322]  = 1;
  ram[5323]  = 1;
  ram[5324]  = 1;
  ram[5325]  = 1;
  ram[5326]  = 1;
  ram[5327]  = 1;
  ram[5328]  = 1;
  ram[5329]  = 1;
  ram[5330]  = 1;
  ram[5331]  = 1;
  ram[5332]  = 1;
  ram[5333]  = 1;
  ram[5334]  = 1;
  ram[5335]  = 1;
  ram[5336]  = 1;
  ram[5337]  = 1;
  ram[5338]  = 1;
  ram[5339]  = 1;
  ram[5340]  = 1;
  ram[5341]  = 1;
  ram[5342]  = 1;
  ram[5343]  = 1;
  ram[5344]  = 1;
  ram[5345]  = 1;
  ram[5346]  = 1;
  ram[5347]  = 1;
  ram[5348]  = 1;
  ram[5349]  = 1;
  ram[5350]  = 1;
  ram[5351]  = 1;
  ram[5352]  = 1;
  ram[5353]  = 1;
  ram[5354]  = 1;
  ram[5355]  = 1;
  ram[5356]  = 1;
  ram[5357]  = 1;
  ram[5358]  = 1;
  ram[5359]  = 1;
  ram[5360]  = 1;
  ram[5361]  = 1;
  ram[5362]  = 1;
  ram[5363]  = 1;
  ram[5364]  = 1;
  ram[5365]  = 1;
  ram[5366]  = 1;
  ram[5367]  = 1;
  ram[5368]  = 1;
  ram[5369]  = 1;
  ram[5370]  = 1;
  ram[5371]  = 1;
  ram[5372]  = 1;
  ram[5373]  = 1;
  ram[5374]  = 1;
  ram[5375]  = 1;
  ram[5376]  = 1;
  ram[5377]  = 1;
  ram[5378]  = 1;
  ram[5379]  = 1;
  ram[5380]  = 1;
  ram[5381]  = 1;
  ram[5382]  = 1;
  ram[5383]  = 1;
  ram[5384]  = 1;
  ram[5385]  = 1;
  ram[5386]  = 1;
  ram[5387]  = 1;
  ram[5388]  = 1;
  ram[5389]  = 1;
  ram[5390]  = 1;
  ram[5391]  = 1;
  ram[5392]  = 1;
  ram[5393]  = 1;
  ram[5394]  = 1;
  ram[5395]  = 1;
  ram[5396]  = 1;
  ram[5397]  = 1;
  ram[5398]  = 1;
  ram[5399]  = 1;
  ram[5400]  = 1;
  ram[5401]  = 1;
  ram[5402]  = 1;
  ram[5403]  = 1;
  ram[5404]  = 1;
  ram[5405]  = 1;
  ram[5406]  = 1;
  ram[5407]  = 1;
  ram[5408]  = 1;
  ram[5409]  = 1;
  ram[5410]  = 1;
  ram[5411]  = 1;
  ram[5412]  = 1;
  ram[5413]  = 1;
  ram[5414]  = 1;
  ram[5415]  = 1;
  ram[5416]  = 1;
  ram[5417]  = 1;
  ram[5418]  = 1;
  ram[5419]  = 1;
  ram[5420]  = 1;
  ram[5421]  = 1;
  ram[5422]  = 1;
  ram[5423]  = 1;
  ram[5424]  = 1;
  ram[5425]  = 1;
  ram[5426]  = 1;
  ram[5427]  = 1;
  ram[5428]  = 1;
  ram[5429]  = 1;
  ram[5430]  = 1;
  ram[5431]  = 1;
  ram[5432]  = 1;
  ram[5433]  = 1;
  ram[5434]  = 1;
  ram[5435]  = 1;
  ram[5436]  = 1;
  ram[5437]  = 1;
  ram[5438]  = 1;
  ram[5439]  = 1;
  ram[5440]  = 1;
  ram[5441]  = 1;
  ram[5442]  = 1;
  ram[5443]  = 1;
  ram[5444]  = 1;
  ram[5445]  = 1;
  ram[5446]  = 1;
  ram[5447]  = 1;
  ram[5448]  = 1;
  ram[5449]  = 1;
  ram[5450]  = 1;
  ram[5451]  = 1;
  ram[5452]  = 1;
  ram[5453]  = 1;
  ram[5454]  = 1;
  ram[5455]  = 1;
  ram[5456]  = 1;
  ram[5457]  = 1;
  ram[5458]  = 1;
  ram[5459]  = 1;
  ram[5460]  = 1;
  ram[5461]  = 1;
  ram[5462]  = 1;
  ram[5463]  = 1;
  ram[5464]  = 1;
  ram[5465]  = 1;
  ram[5466]  = 1;
  ram[5467]  = 1;
  ram[5468]  = 1;
  ram[5469]  = 1;
  ram[5470]  = 1;
  ram[5471]  = 1;
  ram[5472]  = 1;
  ram[5473]  = 1;
  ram[5474]  = 1;
  ram[5475]  = 1;
  ram[5476]  = 1;
  ram[5477]  = 1;
  ram[5478]  = 1;
  ram[5479]  = 1;
  ram[5480]  = 1;
  ram[5481]  = 1;
  ram[5482]  = 1;
  ram[5483]  = 1;
  ram[5484]  = 1;
  ram[5485]  = 1;
  ram[5486]  = 1;
  ram[5487]  = 1;
  ram[5488]  = 1;
  ram[5489]  = 1;
  ram[5490]  = 1;
  ram[5491]  = 1;
  ram[5492]  = 1;
  ram[5493]  = 1;
  ram[5494]  = 1;
  ram[5495]  = 1;
  ram[5496]  = 1;
  ram[5497]  = 1;
  ram[5498]  = 1;
  ram[5499]  = 1;
  ram[5500]  = 1;
  ram[5501]  = 1;
  ram[5502]  = 1;
  ram[5503]  = 1;
  ram[5504]  = 1;
  ram[5505]  = 1;
  ram[5506]  = 1;
  ram[5507]  = 1;
  ram[5508]  = 1;
  ram[5509]  = 1;
  ram[5510]  = 1;
  ram[5511]  = 1;
  ram[5512]  = 1;
  ram[5513]  = 1;
  ram[5514]  = 1;
  ram[5515]  = 1;
  ram[5516]  = 1;
  ram[5517]  = 1;
  ram[5518]  = 1;
  ram[5519]  = 1;
  ram[5520]  = 1;
  ram[5521]  = 1;
  ram[5522]  = 1;
  ram[5523]  = 1;
  ram[5524]  = 1;
  ram[5525]  = 1;
  ram[5526]  = 1;
  ram[5527]  = 1;
  ram[5528]  = 1;
  ram[5529]  = 1;
  ram[5530]  = 1;
  ram[5531]  = 1;
  ram[5532]  = 1;
  ram[5533]  = 1;
  ram[5534]  = 1;
  ram[5535]  = 1;
  ram[5536]  = 1;
  ram[5537]  = 1;
  ram[5538]  = 1;
  ram[5539]  = 1;
  ram[5540]  = 1;
  ram[5541]  = 1;
  ram[5542]  = 1;
  ram[5543]  = 1;
  ram[5544]  = 1;
  ram[5545]  = 1;
  ram[5546]  = 1;
  ram[5547]  = 1;
  ram[5548]  = 1;
  ram[5549]  = 1;
  ram[5550]  = 1;
  ram[5551]  = 1;
  ram[5552]  = 1;
  ram[5553]  = 1;
  ram[5554]  = 1;
  ram[5555]  = 1;
  ram[5556]  = 1;
  ram[5557]  = 1;
  ram[5558]  = 1;
  ram[5559]  = 1;
  ram[5560]  = 1;
  ram[5561]  = 1;
  ram[5562]  = 1;
  ram[5563]  = 1;
  ram[5564]  = 1;
  ram[5565]  = 1;
  ram[5566]  = 1;
  ram[5567]  = 1;
  ram[5568]  = 1;
  ram[5569]  = 1;
  ram[5570]  = 1;
  ram[5571]  = 1;
  ram[5572]  = 1;
  ram[5573]  = 1;
  ram[5574]  = 1;
  ram[5575]  = 1;
  ram[5576]  = 1;
  ram[5577]  = 1;
  ram[5578]  = 1;
  ram[5579]  = 1;
  ram[5580]  = 1;
  ram[5581]  = 1;
  ram[5582]  = 1;
  ram[5583]  = 1;
  ram[5584]  = 1;
  ram[5585]  = 1;
  ram[5586]  = 1;
  ram[5587]  = 1;
  ram[5588]  = 1;
  ram[5589]  = 1;
  ram[5590]  = 1;
  ram[5591]  = 1;
  ram[5592]  = 1;
  ram[5593]  = 1;
  ram[5594]  = 1;
  ram[5595]  = 1;
  ram[5596]  = 1;
  ram[5597]  = 1;
  ram[5598]  = 1;
  ram[5599]  = 1;
  ram[5600]  = 1;
  ram[5601]  = 1;
  ram[5602]  = 1;
  ram[5603]  = 1;
  ram[5604]  = 1;
  ram[5605]  = 1;
  ram[5606]  = 1;
  ram[5607]  = 1;
  ram[5608]  = 1;
  ram[5609]  = 1;
  ram[5610]  = 1;
  ram[5611]  = 1;
  ram[5612]  = 1;
  ram[5613]  = 1;
  ram[5614]  = 1;
  ram[5615]  = 1;
  ram[5616]  = 1;
  ram[5617]  = 1;
  ram[5618]  = 1;
  ram[5619]  = 1;
  ram[5620]  = 1;
  ram[5621]  = 1;
  ram[5622]  = 1;
  ram[5623]  = 1;
  ram[5624]  = 1;
  ram[5625]  = 1;
  ram[5626]  = 1;
  ram[5627]  = 1;
  ram[5628]  = 1;
  ram[5629]  = 1;
  ram[5630]  = 1;
  ram[5631]  = 1;
  ram[5632]  = 1;
  ram[5633]  = 1;
  ram[5634]  = 1;
  ram[5635]  = 1;
  ram[5636]  = 1;
  ram[5637]  = 1;
  ram[5638]  = 1;
  ram[5639]  = 1;
  ram[5640]  = 1;
  ram[5641]  = 1;
  ram[5642]  = 1;
  ram[5643]  = 1;
  ram[5644]  = 1;
  ram[5645]  = 1;
  ram[5646]  = 1;
  ram[5647]  = 1;
  ram[5648]  = 1;
  ram[5649]  = 1;
  ram[5650]  = 1;
  ram[5651]  = 1;
  ram[5652]  = 1;
  ram[5653]  = 1;
  ram[5654]  = 1;
  ram[5655]  = 1;
  ram[5656]  = 1;
  ram[5657]  = 1;
  ram[5658]  = 1;
  ram[5659]  = 1;
  ram[5660]  = 1;
  ram[5661]  = 1;
  ram[5662]  = 1;
  ram[5663]  = 1;
  ram[5664]  = 1;
  ram[5665]  = 1;
  ram[5666]  = 1;
  ram[5667]  = 1;
  ram[5668]  = 1;
  ram[5669]  = 1;
  ram[5670]  = 1;
  ram[5671]  = 1;
  ram[5672]  = 1;
  ram[5673]  = 1;
  ram[5674]  = 1;
  ram[5675]  = 1;
  ram[5676]  = 1;
  ram[5677]  = 1;
  ram[5678]  = 1;
  ram[5679]  = 1;
  ram[5680]  = 1;
  ram[5681]  = 1;
  ram[5682]  = 1;
  ram[5683]  = 1;
  ram[5684]  = 1;
  ram[5685]  = 1;
  ram[5686]  = 1;
  ram[5687]  = 1;
  ram[5688]  = 1;
  ram[5689]  = 1;
  ram[5690]  = 1;
  ram[5691]  = 1;
  ram[5692]  = 1;
  ram[5693]  = 1;
  ram[5694]  = 1;
  ram[5695]  = 1;
  ram[5696]  = 1;
  ram[5697]  = 1;
  ram[5698]  = 1;
  ram[5699]  = 1;
  ram[5700]  = 1;
  ram[5701]  = 1;
  ram[5702]  = 1;
  ram[5703]  = 1;
  ram[5704]  = 1;
  ram[5705]  = 1;
  ram[5706]  = 1;
  ram[5707]  = 1;
  ram[5708]  = 1;
  ram[5709]  = 1;
  ram[5710]  = 1;
  ram[5711]  = 1;
  ram[5712]  = 1;
  ram[5713]  = 1;
  ram[5714]  = 1;
  ram[5715]  = 1;
  ram[5716]  = 1;
  ram[5717]  = 1;
  ram[5718]  = 1;
  ram[5719]  = 1;
  ram[5720]  = 1;
  ram[5721]  = 1;
  ram[5722]  = 1;
  ram[5723]  = 1;
  ram[5724]  = 1;
  ram[5725]  = 1;
  ram[5726]  = 1;
  ram[5727]  = 1;
  ram[5728]  = 1;
  ram[5729]  = 1;
  ram[5730]  = 1;
  ram[5731]  = 1;
  ram[5732]  = 1;
  ram[5733]  = 1;
  ram[5734]  = 1;
  ram[5735]  = 1;
  ram[5736]  = 1;
  ram[5737]  = 1;
  ram[5738]  = 1;
  ram[5739]  = 1;
  ram[5740]  = 1;
  ram[5741]  = 1;
  ram[5742]  = 1;
  ram[5743]  = 1;
  ram[5744]  = 1;
  ram[5745]  = 1;
  ram[5746]  = 1;
  ram[5747]  = 1;
  ram[5748]  = 1;
  ram[5749]  = 1;
  ram[5750]  = 1;
  ram[5751]  = 1;
  ram[5752]  = 1;
  ram[5753]  = 1;
  ram[5754]  = 1;
  ram[5755]  = 1;
  ram[5756]  = 1;
  ram[5757]  = 1;
  ram[5758]  = 1;
  ram[5759]  = 1;
  ram[5760]  = 1;
  ram[5761]  = 1;
  ram[5762]  = 1;
  ram[5763]  = 1;
  ram[5764]  = 1;
  ram[5765]  = 1;
  ram[5766]  = 1;
  ram[5767]  = 1;
  ram[5768]  = 1;
  ram[5769]  = 1;
  ram[5770]  = 1;
  ram[5771]  = 1;
  ram[5772]  = 1;
  ram[5773]  = 1;
  ram[5774]  = 1;
  ram[5775]  = 1;
  ram[5776]  = 1;
  ram[5777]  = 1;
  ram[5778]  = 1;
  ram[5779]  = 1;
  ram[5780]  = 1;
  ram[5781]  = 1;
  ram[5782]  = 1;
  ram[5783]  = 1;
  ram[5784]  = 1;
  ram[5785]  = 1;
  ram[5786]  = 1;
  ram[5787]  = 1;
  ram[5788]  = 1;
  ram[5789]  = 1;
  ram[5790]  = 1;
  ram[5791]  = 1;
  ram[5792]  = 1;
  ram[5793]  = 1;
  ram[5794]  = 1;
  ram[5795]  = 1;
  ram[5796]  = 1;
  ram[5797]  = 1;
  ram[5798]  = 1;
  ram[5799]  = 1;
  ram[5800]  = 1;
  ram[5801]  = 1;
  ram[5802]  = 1;
  ram[5803]  = 1;
  ram[5804]  = 1;
  ram[5805]  = 1;
  ram[5806]  = 1;
  ram[5807]  = 1;
  ram[5808]  = 1;
  ram[5809]  = 1;
  ram[5810]  = 1;
  ram[5811]  = 1;
  ram[5812]  = 1;
  ram[5813]  = 1;
  ram[5814]  = 1;
  ram[5815]  = 1;
  ram[5816]  = 1;
  ram[5817]  = 1;
  ram[5818]  = 1;
  ram[5819]  = 1;
  ram[5820]  = 1;
  ram[5821]  = 1;
  ram[5822]  = 1;
  ram[5823]  = 1;
  ram[5824]  = 1;
  ram[5825]  = 1;
  ram[5826]  = 1;
  ram[5827]  = 1;
  ram[5828]  = 1;
  ram[5829]  = 1;
  ram[5830]  = 1;
  ram[5831]  = 1;
  ram[5832]  = 1;
  ram[5833]  = 1;
  ram[5834]  = 1;
  ram[5835]  = 1;
  ram[5836]  = 1;
  ram[5837]  = 1;
  ram[5838]  = 1;
  ram[5839]  = 1;
  ram[5840]  = 1;
  ram[5841]  = 1;
  ram[5842]  = 1;
  ram[5843]  = 1;
  ram[5844]  = 1;
  ram[5845]  = 1;
  ram[5846]  = 1;
  ram[5847]  = 1;
  ram[5848]  = 1;
  ram[5849]  = 1;
  ram[5850]  = 1;
  ram[5851]  = 1;
  ram[5852]  = 1;
  ram[5853]  = 1;
  ram[5854]  = 1;
  ram[5855]  = 1;
  ram[5856]  = 1;
  ram[5857]  = 1;
  ram[5858]  = 1;
  ram[5859]  = 1;
  ram[5860]  = 1;
  ram[5861]  = 1;
  ram[5862]  = 1;
  ram[5863]  = 1;
  ram[5864]  = 1;
  ram[5865]  = 1;
  ram[5866]  = 1;
  ram[5867]  = 1;
  ram[5868]  = 1;
  ram[5869]  = 1;
  ram[5870]  = 1;
  ram[5871]  = 1;
  ram[5872]  = 1;
  ram[5873]  = 1;
  ram[5874]  = 1;
  ram[5875]  = 1;
  ram[5876]  = 1;
  ram[5877]  = 1;
  ram[5878]  = 1;
  ram[5879]  = 1;
  ram[5880]  = 1;
  ram[5881]  = 1;
  ram[5882]  = 1;
  ram[5883]  = 1;
  ram[5884]  = 1;
  ram[5885]  = 1;
  ram[5886]  = 1;
  ram[5887]  = 1;
  ram[5888]  = 1;
  ram[5889]  = 1;
  ram[5890]  = 1;
  ram[5891]  = 1;
  ram[5892]  = 1;
  ram[5893]  = 1;
  ram[5894]  = 1;
  ram[5895]  = 1;
  ram[5896]  = 1;
  ram[5897]  = 1;
  ram[5898]  = 1;
  ram[5899]  = 1;
  ram[5900]  = 1;
  ram[5901]  = 1;
  ram[5902]  = 1;
  ram[5903]  = 1;
  ram[5904]  = 1;
  ram[5905]  = 1;
  ram[5906]  = 1;
  ram[5907]  = 1;
  ram[5908]  = 1;
  ram[5909]  = 1;
  ram[5910]  = 1;
  ram[5911]  = 1;
  ram[5912]  = 1;
  ram[5913]  = 1;
  ram[5914]  = 1;
  ram[5915]  = 1;
  ram[5916]  = 1;
  ram[5917]  = 1;
  ram[5918]  = 1;
  ram[5919]  = 1;
  ram[5920]  = 1;
  ram[5921]  = 1;
  ram[5922]  = 1;
  ram[5923]  = 1;
  ram[5924]  = 1;
  ram[5925]  = 1;
  ram[5926]  = 1;
  ram[5927]  = 1;
  ram[5928]  = 1;
  ram[5929]  = 1;
  ram[5930]  = 1;
  ram[5931]  = 1;
  ram[5932]  = 1;
  ram[5933]  = 1;
  ram[5934]  = 1;
  ram[5935]  = 1;
  ram[5936]  = 1;
  ram[5937]  = 1;
  ram[5938]  = 1;
  ram[5939]  = 1;
  ram[5940]  = 1;
  ram[5941]  = 1;
  ram[5942]  = 1;
  ram[5943]  = 1;
  ram[5944]  = 1;
  ram[5945]  = 1;
  ram[5946]  = 1;
  ram[5947]  = 1;
  ram[5948]  = 1;
  ram[5949]  = 1;
  ram[5950]  = 1;
  ram[5951]  = 1;
  ram[5952]  = 1;
  ram[5953]  = 1;
  ram[5954]  = 1;
  ram[5955]  = 1;
  ram[5956]  = 1;
  ram[5957]  = 1;
  ram[5958]  = 1;
  ram[5959]  = 1;
  ram[5960]  = 1;
  ram[5961]  = 1;
  ram[5962]  = 1;
  ram[5963]  = 1;
  ram[5964]  = 1;
  ram[5965]  = 1;
  ram[5966]  = 1;
  ram[5967]  = 1;
  ram[5968]  = 1;
  ram[5969]  = 1;
  ram[5970]  = 1;
  ram[5971]  = 1;
  ram[5972]  = 1;
  ram[5973]  = 1;
  ram[5974]  = 1;
  ram[5975]  = 1;
  ram[5976]  = 1;
  ram[5977]  = 1;
  ram[5978]  = 1;
  ram[5979]  = 1;
  ram[5980]  = 1;
  ram[5981]  = 1;
  ram[5982]  = 1;
  ram[5983]  = 1;
  ram[5984]  = 1;
  ram[5985]  = 1;
  ram[5986]  = 1;
  ram[5987]  = 1;
  ram[5988]  = 1;
  ram[5989]  = 1;
  ram[5990]  = 1;
  ram[5991]  = 1;
  ram[5992]  = 1;
  ram[5993]  = 1;
  ram[5994]  = 1;
  ram[5995]  = 1;
  ram[5996]  = 1;
  ram[5997]  = 1;
  ram[5998]  = 1;
  ram[5999]  = 1;
  ram[6000]  = 1;
  ram[6001]  = 1;
  ram[6002]  = 1;
  ram[6003]  = 1;
  ram[6004]  = 1;
  ram[6005]  = 1;
  ram[6006]  = 1;
  ram[6007]  = 1;
  ram[6008]  = 1;
  ram[6009]  = 1;
  ram[6010]  = 1;
  ram[6011]  = 1;
  ram[6012]  = 1;
  ram[6013]  = 1;
  ram[6014]  = 1;
  ram[6015]  = 1;
  ram[6016]  = 1;
  ram[6017]  = 1;
  ram[6018]  = 1;
  ram[6019]  = 1;
  ram[6020]  = 1;
  ram[6021]  = 1;
  ram[6022]  = 1;
  ram[6023]  = 1;
  ram[6024]  = 1;
  ram[6025]  = 1;
  ram[6026]  = 1;
  ram[6027]  = 1;
  ram[6028]  = 1;
  ram[6029]  = 1;
  ram[6030]  = 1;
  ram[6031]  = 1;
  ram[6032]  = 1;
  ram[6033]  = 1;
  ram[6034]  = 1;
  ram[6035]  = 1;
  ram[6036]  = 1;
  ram[6037]  = 1;
  ram[6038]  = 1;
  ram[6039]  = 1;
  ram[6040]  = 1;
  ram[6041]  = 1;
  ram[6042]  = 1;
  ram[6043]  = 0;
  ram[6044]  = 0;
  ram[6045]  = 1;
  ram[6046]  = 1;
  ram[6047]  = 1;
  ram[6048]  = 1;
  ram[6049]  = 1;
  ram[6050]  = 1;
  ram[6051]  = 1;
  ram[6052]  = 1;
  ram[6053]  = 1;
  ram[6054]  = 1;
  ram[6055]  = 1;
  ram[6056]  = 1;
  ram[6057]  = 1;
  ram[6058]  = 1;
  ram[6059]  = 1;
  ram[6060]  = 1;
  ram[6061]  = 1;
  ram[6062]  = 1;
  ram[6063]  = 1;
  ram[6064]  = 1;
  ram[6065]  = 1;
  ram[6066]  = 1;
  ram[6067]  = 1;
  ram[6068]  = 1;
  ram[6069]  = 1;
  ram[6070]  = 1;
  ram[6071]  = 1;
  ram[6072]  = 1;
  ram[6073]  = 1;
  ram[6074]  = 1;
  ram[6075]  = 1;
  ram[6076]  = 1;
  ram[6077]  = 1;
  ram[6078]  = 1;
  ram[6079]  = 1;
  ram[6080]  = 1;
  ram[6081]  = 1;
  ram[6082]  = 1;
  ram[6083]  = 1;
  ram[6084]  = 1;
  ram[6085]  = 1;
  ram[6086]  = 1;
  ram[6087]  = 1;
  ram[6088]  = 1;
  ram[6089]  = 1;
  ram[6090]  = 1;
  ram[6091]  = 1;
  ram[6092]  = 1;
  ram[6093]  = 1;
  ram[6094]  = 1;
  ram[6095]  = 1;
  ram[6096]  = 1;
  ram[6097]  = 1;
  ram[6098]  = 1;
  ram[6099]  = 1;
  ram[6100]  = 1;
  ram[6101]  = 1;
  ram[6102]  = 1;
  ram[6103]  = 1;
  ram[6104]  = 1;
  ram[6105]  = 1;
  ram[6106]  = 1;
  ram[6107]  = 1;
  ram[6108]  = 1;
  ram[6109]  = 1;
  ram[6110]  = 1;
  ram[6111]  = 1;
  ram[6112]  = 1;
  ram[6113]  = 1;
  ram[6114]  = 1;
  ram[6115]  = 1;
  ram[6116]  = 1;
  ram[6117]  = 1;
  ram[6118]  = 1;
  ram[6119]  = 1;
  ram[6120]  = 0;
  ram[6121]  = 1;
  ram[6122]  = 1;
  ram[6123]  = 1;
  ram[6124]  = 1;
  ram[6125]  = 1;
  ram[6126]  = 1;
  ram[6127]  = 1;
  ram[6128]  = 1;
  ram[6129]  = 1;
  ram[6130]  = 1;
  ram[6131]  = 1;
  ram[6132]  = 1;
  ram[6133]  = 1;
  ram[6134]  = 1;
  ram[6135]  = 1;
  ram[6136]  = 0;
  ram[6137]  = 0;
  ram[6138]  = 0;
  ram[6139]  = 1;
  ram[6140]  = 1;
  ram[6141]  = 1;
  ram[6142]  = 1;
  ram[6143]  = 1;
  ram[6144]  = 1;
  ram[6145]  = 1;
  ram[6146]  = 1;
  ram[6147]  = 1;
  ram[6148]  = 1;
  ram[6149]  = 1;
  ram[6150]  = 1;
  ram[6151]  = 1;
  ram[6152]  = 1;
  ram[6153]  = 1;
  ram[6154]  = 1;
  ram[6155]  = 1;
  ram[6156]  = 1;
  ram[6157]  = 1;
  ram[6158]  = 1;
  ram[6159]  = 1;
  ram[6160]  = 1;
  ram[6161]  = 1;
  ram[6162]  = 1;
  ram[6163]  = 1;
  ram[6164]  = 1;
  ram[6165]  = 1;
  ram[6166]  = 1;
  ram[6167]  = 1;
  ram[6168]  = 1;
  ram[6169]  = 1;
  ram[6170]  = 1;
  ram[6171]  = 1;
  ram[6172]  = 1;
  ram[6173]  = 1;
  ram[6174]  = 1;
  ram[6175]  = 1;
  ram[6176]  = 1;
  ram[6177]  = 1;
  ram[6178]  = 1;
  ram[6179]  = 1;
  ram[6180]  = 1;
  ram[6181]  = 1;
  ram[6182]  = 1;
  ram[6183]  = 1;
  ram[6184]  = 1;
  ram[6185]  = 1;
  ram[6186]  = 1;
  ram[6187]  = 1;
  ram[6188]  = 1;
  ram[6189]  = 1;
  ram[6190]  = 1;
  ram[6191]  = 1;
  ram[6192]  = 1;
  ram[6193]  = 1;
  ram[6194]  = 1;
  ram[6195]  = 1;
  ram[6196]  = 1;
  ram[6197]  = 1;
  ram[6198]  = 1;
  ram[6199]  = 1;
  ram[6200]  = 1;
  ram[6201]  = 1;
  ram[6202]  = 1;
  ram[6203]  = 1;
  ram[6204]  = 1;
  ram[6205]  = 1;
  ram[6206]  = 1;
  ram[6207]  = 1;
  ram[6208]  = 1;
  ram[6209]  = 1;
  ram[6210]  = 1;
  ram[6211]  = 1;
  ram[6212]  = 1;
  ram[6213]  = 1;
  ram[6214]  = 1;
  ram[6215]  = 1;
  ram[6216]  = 1;
  ram[6217]  = 1;
  ram[6218]  = 1;
  ram[6219]  = 1;
  ram[6220]  = 1;
  ram[6221]  = 1;
  ram[6222]  = 1;
  ram[6223]  = 1;
  ram[6224]  = 1;
  ram[6225]  = 1;
  ram[6226]  = 1;
  ram[6227]  = 1;
  ram[6228]  = 1;
  ram[6229]  = 1;
  ram[6230]  = 1;
  ram[6231]  = 1;
  ram[6232]  = 1;
  ram[6233]  = 1;
  ram[6234]  = 1;
  ram[6235]  = 1;
  ram[6236]  = 1;
  ram[6237]  = 1;
  ram[6238]  = 1;
  ram[6239]  = 1;
  ram[6240]  = 1;
  ram[6241]  = 1;
  ram[6242]  = 1;
  ram[6243]  = 0;
  ram[6244]  = 0;
  ram[6245]  = 1;
  ram[6246]  = 1;
  ram[6247]  = 1;
  ram[6248]  = 1;
  ram[6249]  = 1;
  ram[6250]  = 1;
  ram[6251]  = 1;
  ram[6252]  = 1;
  ram[6253]  = 1;
  ram[6254]  = 1;
  ram[6255]  = 1;
  ram[6256]  = 1;
  ram[6257]  = 1;
  ram[6258]  = 1;
  ram[6259]  = 1;
  ram[6260]  = 1;
  ram[6261]  = 1;
  ram[6262]  = 1;
  ram[6263]  = 1;
  ram[6264]  = 1;
  ram[6265]  = 1;
  ram[6266]  = 1;
  ram[6267]  = 1;
  ram[6268]  = 1;
  ram[6269]  = 1;
  ram[6270]  = 1;
  ram[6271]  = 1;
  ram[6272]  = 1;
  ram[6273]  = 1;
  ram[6274]  = 1;
  ram[6275]  = 1;
  ram[6276]  = 1;
  ram[6277]  = 1;
  ram[6278]  = 1;
  ram[6279]  = 1;
  ram[6280]  = 1;
  ram[6281]  = 0;
  ram[6282]  = 0;
  ram[6283]  = 1;
  ram[6284]  = 1;
  ram[6285]  = 1;
  ram[6286]  = 1;
  ram[6287]  = 1;
  ram[6288]  = 1;
  ram[6289]  = 1;
  ram[6290]  = 1;
  ram[6291]  = 1;
  ram[6292]  = 1;
  ram[6293]  = 1;
  ram[6294]  = 1;
  ram[6295]  = 1;
  ram[6296]  = 1;
  ram[6297]  = 1;
  ram[6298]  = 1;
  ram[6299]  = 1;
  ram[6300]  = 1;
  ram[6301]  = 1;
  ram[6302]  = 1;
  ram[6303]  = 1;
  ram[6304]  = 1;
  ram[6305]  = 1;
  ram[6306]  = 1;
  ram[6307]  = 1;
  ram[6308]  = 1;
  ram[6309]  = 1;
  ram[6310]  = 1;
  ram[6311]  = 1;
  ram[6312]  = 1;
  ram[6313]  = 1;
  ram[6314]  = 1;
  ram[6315]  = 1;
  ram[6316]  = 1;
  ram[6317]  = 1;
  ram[6318]  = 1;
  ram[6319]  = 0;
  ram[6320]  = 0;
  ram[6321]  = 1;
  ram[6322]  = 1;
  ram[6323]  = 1;
  ram[6324]  = 1;
  ram[6325]  = 1;
  ram[6326]  = 1;
  ram[6327]  = 1;
  ram[6328]  = 1;
  ram[6329]  = 1;
  ram[6330]  = 1;
  ram[6331]  = 1;
  ram[6332]  = 1;
  ram[6333]  = 1;
  ram[6334]  = 1;
  ram[6335]  = 1;
  ram[6336]  = 0;
  ram[6337]  = 0;
  ram[6338]  = 0;
  ram[6339]  = 0;
  ram[6340]  = 1;
  ram[6341]  = 1;
  ram[6342]  = 1;
  ram[6343]  = 1;
  ram[6344]  = 1;
  ram[6345]  = 1;
  ram[6346]  = 1;
  ram[6347]  = 1;
  ram[6348]  = 1;
  ram[6349]  = 1;
  ram[6350]  = 1;
  ram[6351]  = 1;
  ram[6352]  = 1;
  ram[6353]  = 1;
  ram[6354]  = 1;
  ram[6355]  = 1;
  ram[6356]  = 1;
  ram[6357]  = 1;
  ram[6358]  = 1;
  ram[6359]  = 1;
  ram[6360]  = 1;
  ram[6361]  = 1;
  ram[6362]  = 1;
  ram[6363]  = 1;
  ram[6364]  = 1;
  ram[6365]  = 1;
  ram[6366]  = 1;
  ram[6367]  = 1;
  ram[6368]  = 1;
  ram[6369]  = 1;
  ram[6370]  = 1;
  ram[6371]  = 1;
  ram[6372]  = 1;
  ram[6373]  = 1;
  ram[6374]  = 1;
  ram[6375]  = 1;
  ram[6376]  = 1;
  ram[6377]  = 1;
  ram[6378]  = 1;
  ram[6379]  = 1;
  ram[6380]  = 1;
  ram[6381]  = 1;
  ram[6382]  = 1;
  ram[6383]  = 1;
  ram[6384]  = 1;
  ram[6385]  = 1;
  ram[6386]  = 1;
  ram[6387]  = 1;
  ram[6388]  = 1;
  ram[6389]  = 1;
  ram[6390]  = 1;
  ram[6391]  = 1;
  ram[6392]  = 1;
  ram[6393]  = 1;
  ram[6394]  = 1;
  ram[6395]  = 1;
  ram[6396]  = 1;
  ram[6397]  = 1;
  ram[6398]  = 1;
  ram[6399]  = 1;
  ram[6400]  = 1;
  ram[6401]  = 1;
  ram[6402]  = 1;
  ram[6403]  = 1;
  ram[6404]  = 1;
  ram[6405]  = 1;
  ram[6406]  = 1;
  ram[6407]  = 1;
  ram[6408]  = 1;
  ram[6409]  = 1;
  ram[6410]  = 1;
  ram[6411]  = 1;
  ram[6412]  = 1;
  ram[6413]  = 1;
  ram[6414]  = 1;
  ram[6415]  = 1;
  ram[6416]  = 1;
  ram[6417]  = 1;
  ram[6418]  = 1;
  ram[6419]  = 1;
  ram[6420]  = 1;
  ram[6421]  = 1;
  ram[6422]  = 1;
  ram[6423]  = 1;
  ram[6424]  = 1;
  ram[6425]  = 1;
  ram[6426]  = 1;
  ram[6427]  = 1;
  ram[6428]  = 1;
  ram[6429]  = 1;
  ram[6430]  = 1;
  ram[6431]  = 1;
  ram[6432]  = 1;
  ram[6433]  = 1;
  ram[6434]  = 1;
  ram[6435]  = 1;
  ram[6436]  = 1;
  ram[6437]  = 1;
  ram[6438]  = 0;
  ram[6439]  = 0;
  ram[6440]  = 1;
  ram[6441]  = 1;
  ram[6442]  = 1;
  ram[6443]  = 0;
  ram[6444]  = 0;
  ram[6445]  = 1;
  ram[6446]  = 1;
  ram[6447]  = 1;
  ram[6448]  = 0;
  ram[6449]  = 1;
  ram[6450]  = 1;
  ram[6451]  = 1;
  ram[6452]  = 1;
  ram[6453]  = 1;
  ram[6454]  = 1;
  ram[6455]  = 1;
  ram[6456]  = 1;
  ram[6457]  = 1;
  ram[6458]  = 1;
  ram[6459]  = 1;
  ram[6460]  = 1;
  ram[6461]  = 1;
  ram[6462]  = 1;
  ram[6463]  = 1;
  ram[6464]  = 1;
  ram[6465]  = 1;
  ram[6466]  = 1;
  ram[6467]  = 1;
  ram[6468]  = 0;
  ram[6469]  = 0;
  ram[6470]  = 0;
  ram[6471]  = 0;
  ram[6472]  = 0;
  ram[6473]  = 0;
  ram[6474]  = 0;
  ram[6475]  = 0;
  ram[6476]  = 0;
  ram[6477]  = 0;
  ram[6478]  = 0;
  ram[6479]  = 1;
  ram[6480]  = 1;
  ram[6481]  = 0;
  ram[6482]  = 0;
  ram[6483]  = 1;
  ram[6484]  = 1;
  ram[6485]  = 1;
  ram[6486]  = 1;
  ram[6487]  = 1;
  ram[6488]  = 1;
  ram[6489]  = 1;
  ram[6490]  = 1;
  ram[6491]  = 1;
  ram[6492]  = 1;
  ram[6493]  = 1;
  ram[6494]  = 1;
  ram[6495]  = 1;
  ram[6496]  = 1;
  ram[6497]  = 1;
  ram[6498]  = 1;
  ram[6499]  = 1;
  ram[6500]  = 1;
  ram[6501]  = 1;
  ram[6502]  = 1;
  ram[6503]  = 1;
  ram[6504]  = 1;
  ram[6505]  = 1;
  ram[6506]  = 1;
  ram[6507]  = 1;
  ram[6508]  = 1;
  ram[6509]  = 1;
  ram[6510]  = 1;
  ram[6511]  = 1;
  ram[6512]  = 1;
  ram[6513]  = 1;
  ram[6514]  = 1;
  ram[6515]  = 1;
  ram[6516]  = 1;
  ram[6517]  = 1;
  ram[6518]  = 1;
  ram[6519]  = 0;
  ram[6520]  = 0;
  ram[6521]  = 1;
  ram[6522]  = 1;
  ram[6523]  = 1;
  ram[6524]  = 1;
  ram[6525]  = 1;
  ram[6526]  = 1;
  ram[6527]  = 1;
  ram[6528]  = 1;
  ram[6529]  = 1;
  ram[6530]  = 1;
  ram[6531]  = 1;
  ram[6532]  = 1;
  ram[6533]  = 1;
  ram[6534]  = 1;
  ram[6535]  = 0;
  ram[6536]  = 0;
  ram[6537]  = 1;
  ram[6538]  = 1;
  ram[6539]  = 0;
  ram[6540]  = 0;
  ram[6541]  = 1;
  ram[6542]  = 1;
  ram[6543]  = 1;
  ram[6544]  = 1;
  ram[6545]  = 1;
  ram[6546]  = 1;
  ram[6547]  = 1;
  ram[6548]  = 1;
  ram[6549]  = 1;
  ram[6550]  = 1;
  ram[6551]  = 1;
  ram[6552]  = 1;
  ram[6553]  = 0;
  ram[6554]  = 0;
  ram[6555]  = 0;
  ram[6556]  = 0;
  ram[6557]  = 0;
  ram[6558]  = 0;
  ram[6559]  = 0;
  ram[6560]  = 0;
  ram[6561]  = 0;
  ram[6562]  = 0;
  ram[6563]  = 0;
  ram[6564]  = 0;
  ram[6565]  = 0;
  ram[6566]  = 0;
  ram[6567]  = 0;
  ram[6568]  = 0;
  ram[6569]  = 0;
  ram[6570]  = 0;
  ram[6571]  = 0;
  ram[6572]  = 0;
  ram[6573]  = 0;
  ram[6574]  = 0;
  ram[6575]  = 0;
  ram[6576]  = 0;
  ram[6577]  = 0;
  ram[6578]  = 0;
  ram[6579]  = 0;
  ram[6580]  = 0;
  ram[6581]  = 0;
  ram[6582]  = 0;
  ram[6583]  = 0;
  ram[6584]  = 1;
  ram[6585]  = 1;
  ram[6586]  = 1;
  ram[6587]  = 1;
  ram[6588]  = 1;
  ram[6589]  = 1;
  ram[6590]  = 1;
  ram[6591]  = 1;
  ram[6592]  = 1;
  ram[6593]  = 1;
  ram[6594]  = 1;
  ram[6595]  = 1;
  ram[6596]  = 1;
  ram[6597]  = 1;
  ram[6598]  = 1;
  ram[6599]  = 1;
  ram[6600]  = 1;
  ram[6601]  = 1;
  ram[6602]  = 1;
  ram[6603]  = 1;
  ram[6604]  = 1;
  ram[6605]  = 1;
  ram[6606]  = 1;
  ram[6607]  = 1;
  ram[6608]  = 1;
  ram[6609]  = 1;
  ram[6610]  = 1;
  ram[6611]  = 1;
  ram[6612]  = 1;
  ram[6613]  = 1;
  ram[6614]  = 1;
  ram[6615]  = 1;
  ram[6616]  = 1;
  ram[6617]  = 1;
  ram[6618]  = 1;
  ram[6619]  = 1;
  ram[6620]  = 1;
  ram[6621]  = 1;
  ram[6622]  = 1;
  ram[6623]  = 1;
  ram[6624]  = 1;
  ram[6625]  = 1;
  ram[6626]  = 1;
  ram[6627]  = 1;
  ram[6628]  = 1;
  ram[6629]  = 1;
  ram[6630]  = 1;
  ram[6631]  = 1;
  ram[6632]  = 1;
  ram[6633]  = 0;
  ram[6634]  = 0;
  ram[6635]  = 0;
  ram[6636]  = 0;
  ram[6637]  = 0;
  ram[6638]  = 0;
  ram[6639]  = 0;
  ram[6640]  = 0;
  ram[6641]  = 1;
  ram[6642]  = 1;
  ram[6643]  = 0;
  ram[6644]  = 0;
  ram[6645]  = 1;
  ram[6646]  = 1;
  ram[6647]  = 0;
  ram[6648]  = 0;
  ram[6649]  = 0;
  ram[6650]  = 1;
  ram[6651]  = 1;
  ram[6652]  = 1;
  ram[6653]  = 1;
  ram[6654]  = 1;
  ram[6655]  = 1;
  ram[6656]  = 1;
  ram[6657]  = 1;
  ram[6658]  = 1;
  ram[6659]  = 1;
  ram[6660]  = 1;
  ram[6661]  = 1;
  ram[6662]  = 1;
  ram[6663]  = 1;
  ram[6664]  = 1;
  ram[6665]  = 1;
  ram[6666]  = 1;
  ram[6667]  = 1;
  ram[6668]  = 0;
  ram[6669]  = 0;
  ram[6670]  = 0;
  ram[6671]  = 0;
  ram[6672]  = 0;
  ram[6673]  = 0;
  ram[6674]  = 0;
  ram[6675]  = 0;
  ram[6676]  = 0;
  ram[6677]  = 0;
  ram[6678]  = 0;
  ram[6679]  = 1;
  ram[6680]  = 1;
  ram[6681]  = 0;
  ram[6682]  = 0;
  ram[6683]  = 1;
  ram[6684]  = 1;
  ram[6685]  = 1;
  ram[6686]  = 1;
  ram[6687]  = 1;
  ram[6688]  = 1;
  ram[6689]  = 1;
  ram[6690]  = 1;
  ram[6691]  = 1;
  ram[6692]  = 1;
  ram[6693]  = 1;
  ram[6694]  = 1;
  ram[6695]  = 1;
  ram[6696]  = 1;
  ram[6697]  = 1;
  ram[6698]  = 1;
  ram[6699]  = 1;
  ram[6700]  = 1;
  ram[6701]  = 1;
  ram[6702]  = 1;
  ram[6703]  = 1;
  ram[6704]  = 1;
  ram[6705]  = 1;
  ram[6706]  = 1;
  ram[6707]  = 1;
  ram[6708]  = 1;
  ram[6709]  = 1;
  ram[6710]  = 1;
  ram[6711]  = 1;
  ram[6712]  = 1;
  ram[6713]  = 1;
  ram[6714]  = 1;
  ram[6715]  = 1;
  ram[6716]  = 1;
  ram[6717]  = 1;
  ram[6718]  = 1;
  ram[6719]  = 0;
  ram[6720]  = 0;
  ram[6721]  = 1;
  ram[6722]  = 1;
  ram[6723]  = 1;
  ram[6724]  = 1;
  ram[6725]  = 1;
  ram[6726]  = 1;
  ram[6727]  = 1;
  ram[6728]  = 1;
  ram[6729]  = 1;
  ram[6730]  = 1;
  ram[6731]  = 1;
  ram[6732]  = 1;
  ram[6733]  = 1;
  ram[6734]  = 0;
  ram[6735]  = 0;
  ram[6736]  = 0;
  ram[6737]  = 1;
  ram[6738]  = 1;
  ram[6739]  = 0;
  ram[6740]  = 0;
  ram[6741]  = 0;
  ram[6742]  = 1;
  ram[6743]  = 1;
  ram[6744]  = 1;
  ram[6745]  = 1;
  ram[6746]  = 1;
  ram[6747]  = 1;
  ram[6748]  = 1;
  ram[6749]  = 1;
  ram[6750]  = 1;
  ram[6751]  = 1;
  ram[6752]  = 1;
  ram[6753]  = 0;
  ram[6754]  = 0;
  ram[6755]  = 0;
  ram[6756]  = 0;
  ram[6757]  = 0;
  ram[6758]  = 0;
  ram[6759]  = 0;
  ram[6760]  = 0;
  ram[6761]  = 0;
  ram[6762]  = 0;
  ram[6763]  = 0;
  ram[6764]  = 0;
  ram[6765]  = 0;
  ram[6766]  = 0;
  ram[6767]  = 0;
  ram[6768]  = 0;
  ram[6769]  = 0;
  ram[6770]  = 0;
  ram[6771]  = 0;
  ram[6772]  = 0;
  ram[6773]  = 0;
  ram[6774]  = 0;
  ram[6775]  = 0;
  ram[6776]  = 0;
  ram[6777]  = 0;
  ram[6778]  = 0;
  ram[6779]  = 0;
  ram[6780]  = 0;
  ram[6781]  = 0;
  ram[6782]  = 0;
  ram[6783]  = 0;
  ram[6784]  = 1;
  ram[6785]  = 1;
  ram[6786]  = 1;
  ram[6787]  = 1;
  ram[6788]  = 1;
  ram[6789]  = 1;
  ram[6790]  = 1;
  ram[6791]  = 1;
  ram[6792]  = 1;
  ram[6793]  = 1;
  ram[6794]  = 1;
  ram[6795]  = 1;
  ram[6796]  = 1;
  ram[6797]  = 1;
  ram[6798]  = 1;
  ram[6799]  = 1;
  ram[6800]  = 1;
  ram[6801]  = 1;
  ram[6802]  = 1;
  ram[6803]  = 1;
  ram[6804]  = 1;
  ram[6805]  = 1;
  ram[6806]  = 1;
  ram[6807]  = 1;
  ram[6808]  = 1;
  ram[6809]  = 1;
  ram[6810]  = 1;
  ram[6811]  = 1;
  ram[6812]  = 1;
  ram[6813]  = 1;
  ram[6814]  = 1;
  ram[6815]  = 1;
  ram[6816]  = 1;
  ram[6817]  = 1;
  ram[6818]  = 1;
  ram[6819]  = 1;
  ram[6820]  = 0;
  ram[6821]  = 0;
  ram[6822]  = 0;
  ram[6823]  = 0;
  ram[6824]  = 0;
  ram[6825]  = 0;
  ram[6826]  = 0;
  ram[6827]  = 0;
  ram[6828]  = 1;
  ram[6829]  = 1;
  ram[6830]  = 0;
  ram[6831]  = 0;
  ram[6832]  = 0;
  ram[6833]  = 0;
  ram[6834]  = 0;
  ram[6835]  = 0;
  ram[6836]  = 0;
  ram[6837]  = 0;
  ram[6838]  = 1;
  ram[6839]  = 1;
  ram[6840]  = 1;
  ram[6841]  = 1;
  ram[6842]  = 1;
  ram[6843]  = 0;
  ram[6844]  = 0;
  ram[6845]  = 1;
  ram[6846]  = 1;
  ram[6847]  = 1;
  ram[6848]  = 0;
  ram[6849]  = 0;
  ram[6850]  = 0;
  ram[6851]  = 1;
  ram[6852]  = 1;
  ram[6853]  = 1;
  ram[6854]  = 1;
  ram[6855]  = 1;
  ram[6856]  = 1;
  ram[6857]  = 0;
  ram[6858]  = 0;
  ram[6859]  = 0;
  ram[6860]  = 0;
  ram[6861]  = 0;
  ram[6862]  = 0;
  ram[6863]  = 0;
  ram[6864]  = 0;
  ram[6865]  = 0;
  ram[6866]  = 1;
  ram[6867]  = 1;
  ram[6868]  = 1;
  ram[6869]  = 1;
  ram[6870]  = 1;
  ram[6871]  = 1;
  ram[6872]  = 1;
  ram[6873]  = 1;
  ram[6874]  = 1;
  ram[6875]  = 1;
  ram[6876]  = 1;
  ram[6877]  = 0;
  ram[6878]  = 0;
  ram[6879]  = 1;
  ram[6880]  = 1;
  ram[6881]  = 0;
  ram[6882]  = 0;
  ram[6883]  = 1;
  ram[6884]  = 1;
  ram[6885]  = 1;
  ram[6886]  = 1;
  ram[6887]  = 1;
  ram[6888]  = 1;
  ram[6889]  = 1;
  ram[6890]  = 1;
  ram[6891]  = 1;
  ram[6892]  = 1;
  ram[6893]  = 1;
  ram[6894]  = 1;
  ram[6895]  = 1;
  ram[6896]  = 1;
  ram[6897]  = 1;
  ram[6898]  = 1;
  ram[6899]  = 1;
  ram[6900]  = 1;
  ram[6901]  = 1;
  ram[6902]  = 1;
  ram[6903]  = 1;
  ram[6904]  = 1;
  ram[6905]  = 1;
  ram[6906]  = 1;
  ram[6907]  = 1;
  ram[6908]  = 1;
  ram[6909]  = 1;
  ram[6910]  = 1;
  ram[6911]  = 1;
  ram[6912]  = 1;
  ram[6913]  = 1;
  ram[6914]  = 1;
  ram[6915]  = 1;
  ram[6916]  = 1;
  ram[6917]  = 1;
  ram[6918]  = 1;
  ram[6919]  = 0;
  ram[6920]  = 1;
  ram[6921]  = 1;
  ram[6922]  = 1;
  ram[6923]  = 1;
  ram[6924]  = 1;
  ram[6925]  = 1;
  ram[6926]  = 1;
  ram[6927]  = 1;
  ram[6928]  = 1;
  ram[6929]  = 1;
  ram[6930]  = 1;
  ram[6931]  = 1;
  ram[6932]  = 1;
  ram[6933]  = 0;
  ram[6934]  = 0;
  ram[6935]  = 0;
  ram[6936]  = 1;
  ram[6937]  = 1;
  ram[6938]  = 1;
  ram[6939]  = 1;
  ram[6940]  = 0;
  ram[6941]  = 0;
  ram[6942]  = 0;
  ram[6943]  = 1;
  ram[6944]  = 1;
  ram[6945]  = 1;
  ram[6946]  = 1;
  ram[6947]  = 1;
  ram[6948]  = 1;
  ram[6949]  = 1;
  ram[6950]  = 1;
  ram[6951]  = 1;
  ram[6952]  = 1;
  ram[6953]  = 0;
  ram[6954]  = 0;
  ram[6955]  = 0;
  ram[6956]  = 0;
  ram[6957]  = 0;
  ram[6958]  = 0;
  ram[6959]  = 0;
  ram[6960]  = 0;
  ram[6961]  = 0;
  ram[6962]  = 0;
  ram[6963]  = 0;
  ram[6964]  = 0;
  ram[6965]  = 0;
  ram[6966]  = 0;
  ram[6967]  = 0;
  ram[6968]  = 0;
  ram[6969]  = 0;
  ram[6970]  = 0;
  ram[6971]  = 0;
  ram[6972]  = 0;
  ram[6973]  = 0;
  ram[6974]  = 0;
  ram[6975]  = 0;
  ram[6976]  = 0;
  ram[6977]  = 0;
  ram[6978]  = 0;
  ram[6979]  = 0;
  ram[6980]  = 0;
  ram[6981]  = 0;
  ram[6982]  = 0;
  ram[6983]  = 0;
  ram[6984]  = 1;
  ram[6985]  = 1;
  ram[6986]  = 1;
  ram[6987]  = 1;
  ram[6988]  = 1;
  ram[6989]  = 1;
  ram[6990]  = 1;
  ram[6991]  = 1;
  ram[6992]  = 1;
  ram[6993]  = 1;
  ram[6994]  = 1;
  ram[6995]  = 1;
  ram[6996]  = 1;
  ram[6997]  = 1;
  ram[6998]  = 1;
  ram[6999]  = 1;
  ram[7000]  = 1;
  ram[7001]  = 1;
  ram[7002]  = 1;
  ram[7003]  = 1;
  ram[7004]  = 1;
  ram[7005]  = 1;
  ram[7006]  = 1;
  ram[7007]  = 1;
  ram[7008]  = 1;
  ram[7009]  = 1;
  ram[7010]  = 1;
  ram[7011]  = 1;
  ram[7012]  = 1;
  ram[7013]  = 1;
  ram[7014]  = 1;
  ram[7015]  = 1;
  ram[7016]  = 1;
  ram[7017]  = 1;
  ram[7018]  = 1;
  ram[7019]  = 1;
  ram[7020]  = 0;
  ram[7021]  = 0;
  ram[7022]  = 1;
  ram[7023]  = 1;
  ram[7024]  = 1;
  ram[7025]  = 1;
  ram[7026]  = 0;
  ram[7027]  = 0;
  ram[7028]  = 1;
  ram[7029]  = 1;
  ram[7030]  = 0;
  ram[7031]  = 0;
  ram[7032]  = 1;
  ram[7033]  = 1;
  ram[7034]  = 0;
  ram[7035]  = 0;
  ram[7036]  = 1;
  ram[7037]  = 1;
  ram[7038]  = 1;
  ram[7039]  = 1;
  ram[7040]  = 1;
  ram[7041]  = 1;
  ram[7042]  = 1;
  ram[7043]  = 0;
  ram[7044]  = 0;
  ram[7045]  = 1;
  ram[7046]  = 1;
  ram[7047]  = 1;
  ram[7048]  = 1;
  ram[7049]  = 1;
  ram[7050]  = 0;
  ram[7051]  = 0;
  ram[7052]  = 1;
  ram[7053]  = 1;
  ram[7054]  = 1;
  ram[7055]  = 1;
  ram[7056]  = 1;
  ram[7057]  = 0;
  ram[7058]  = 0;
  ram[7059]  = 0;
  ram[7060]  = 1;
  ram[7061]  = 1;
  ram[7062]  = 1;
  ram[7063]  = 0;
  ram[7064]  = 0;
  ram[7065]  = 0;
  ram[7066]  = 1;
  ram[7067]  = 1;
  ram[7068]  = 1;
  ram[7069]  = 1;
  ram[7070]  = 1;
  ram[7071]  = 1;
  ram[7072]  = 1;
  ram[7073]  = 1;
  ram[7074]  = 1;
  ram[7075]  = 1;
  ram[7076]  = 0;
  ram[7077]  = 0;
  ram[7078]  = 0;
  ram[7079]  = 1;
  ram[7080]  = 1;
  ram[7081]  = 0;
  ram[7082]  = 0;
  ram[7083]  = 1;
  ram[7084]  = 1;
  ram[7085]  = 1;
  ram[7086]  = 1;
  ram[7087]  = 1;
  ram[7088]  = 1;
  ram[7089]  = 1;
  ram[7090]  = 1;
  ram[7091]  = 1;
  ram[7092]  = 1;
  ram[7093]  = 1;
  ram[7094]  = 1;
  ram[7095]  = 1;
  ram[7096]  = 1;
  ram[7097]  = 1;
  ram[7098]  = 1;
  ram[7099]  = 1;
  ram[7100]  = 1;
  ram[7101]  = 1;
  ram[7102]  = 1;
  ram[7103]  = 1;
  ram[7104]  = 1;
  ram[7105]  = 1;
  ram[7106]  = 1;
  ram[7107]  = 1;
  ram[7108]  = 1;
  ram[7109]  = 1;
  ram[7110]  = 1;
  ram[7111]  = 1;
  ram[7112]  = 1;
  ram[7113]  = 1;
  ram[7114]  = 1;
  ram[7115]  = 0;
  ram[7116]  = 0;
  ram[7117]  = 0;
  ram[7118]  = 0;
  ram[7119]  = 0;
  ram[7120]  = 0;
  ram[7121]  = 0;
  ram[7122]  = 0;
  ram[7123]  = 0;
  ram[7124]  = 0;
  ram[7125]  = 0;
  ram[7126]  = 0;
  ram[7127]  = 1;
  ram[7128]  = 1;
  ram[7129]  = 1;
  ram[7130]  = 1;
  ram[7131]  = 1;
  ram[7132]  = 0;
  ram[7133]  = 0;
  ram[7134]  = 0;
  ram[7135]  = 1;
  ram[7136]  = 1;
  ram[7137]  = 1;
  ram[7138]  = 1;
  ram[7139]  = 1;
  ram[7140]  = 1;
  ram[7141]  = 0;
  ram[7142]  = 0;
  ram[7143]  = 0;
  ram[7144]  = 1;
  ram[7145]  = 1;
  ram[7146]  = 1;
  ram[7147]  = 1;
  ram[7148]  = 1;
  ram[7149]  = 1;
  ram[7150]  = 1;
  ram[7151]  = 1;
  ram[7152]  = 1;
  ram[7153]  = 1;
  ram[7154]  = 1;
  ram[7155]  = 1;
  ram[7156]  = 1;
  ram[7157]  = 1;
  ram[7158]  = 1;
  ram[7159]  = 1;
  ram[7160]  = 1;
  ram[7161]  = 1;
  ram[7162]  = 1;
  ram[7163]  = 1;
  ram[7164]  = 1;
  ram[7165]  = 1;
  ram[7166]  = 1;
  ram[7167]  = 1;
  ram[7168]  = 1;
  ram[7169]  = 1;
  ram[7170]  = 1;
  ram[7171]  = 1;
  ram[7172]  = 1;
  ram[7173]  = 1;
  ram[7174]  = 1;
  ram[7175]  = 1;
  ram[7176]  = 1;
  ram[7177]  = 1;
  ram[7178]  = 1;
  ram[7179]  = 1;
  ram[7180]  = 0;
  ram[7181]  = 0;
  ram[7182]  = 0;
  ram[7183]  = 0;
  ram[7184]  = 1;
  ram[7185]  = 1;
  ram[7186]  = 1;
  ram[7187]  = 1;
  ram[7188]  = 1;
  ram[7189]  = 1;
  ram[7190]  = 1;
  ram[7191]  = 1;
  ram[7192]  = 1;
  ram[7193]  = 1;
  ram[7194]  = 1;
  ram[7195]  = 1;
  ram[7196]  = 1;
  ram[7197]  = 1;
  ram[7198]  = 1;
  ram[7199]  = 1;
  ram[7200]  = 1;
  ram[7201]  = 1;
  ram[7202]  = 1;
  ram[7203]  = 1;
  ram[7204]  = 1;
  ram[7205]  = 1;
  ram[7206]  = 1;
  ram[7207]  = 1;
  ram[7208]  = 1;
  ram[7209]  = 1;
  ram[7210]  = 1;
  ram[7211]  = 1;
  ram[7212]  = 1;
  ram[7213]  = 1;
  ram[7214]  = 1;
  ram[7215]  = 1;
  ram[7216]  = 1;
  ram[7217]  = 1;
  ram[7218]  = 1;
  ram[7219]  = 1;
  ram[7220]  = 0;
  ram[7221]  = 0;
  ram[7222]  = 1;
  ram[7223]  = 1;
  ram[7224]  = 1;
  ram[7225]  = 1;
  ram[7226]  = 0;
  ram[7227]  = 0;
  ram[7228]  = 1;
  ram[7229]  = 1;
  ram[7230]  = 1;
  ram[7231]  = 1;
  ram[7232]  = 1;
  ram[7233]  = 1;
  ram[7234]  = 1;
  ram[7235]  = 0;
  ram[7236]  = 1;
  ram[7237]  = 1;
  ram[7238]  = 1;
  ram[7239]  = 1;
  ram[7240]  = 1;
  ram[7241]  = 1;
  ram[7242]  = 1;
  ram[7243]  = 0;
  ram[7244]  = 0;
  ram[7245]  = 1;
  ram[7246]  = 1;
  ram[7247]  = 1;
  ram[7248]  = 1;
  ram[7249]  = 1;
  ram[7250]  = 0;
  ram[7251]  = 0;
  ram[7252]  = 1;
  ram[7253]  = 1;
  ram[7254]  = 1;
  ram[7255]  = 1;
  ram[7256]  = 1;
  ram[7257]  = 0;
  ram[7258]  = 0;
  ram[7259]  = 1;
  ram[7260]  = 1;
  ram[7261]  = 1;
  ram[7262]  = 1;
  ram[7263]  = 1;
  ram[7264]  = 0;
  ram[7265]  = 0;
  ram[7266]  = 1;
  ram[7267]  = 1;
  ram[7268]  = 1;
  ram[7269]  = 1;
  ram[7270]  = 1;
  ram[7271]  = 1;
  ram[7272]  = 1;
  ram[7273]  = 1;
  ram[7274]  = 1;
  ram[7275]  = 1;
  ram[7276]  = 0;
  ram[7277]  = 0;
  ram[7278]  = 1;
  ram[7279]  = 1;
  ram[7280]  = 1;
  ram[7281]  = 0;
  ram[7282]  = 0;
  ram[7283]  = 1;
  ram[7284]  = 1;
  ram[7285]  = 1;
  ram[7286]  = 1;
  ram[7287]  = 1;
  ram[7288]  = 1;
  ram[7289]  = 1;
  ram[7290]  = 1;
  ram[7291]  = 1;
  ram[7292]  = 1;
  ram[7293]  = 1;
  ram[7294]  = 1;
  ram[7295]  = 1;
  ram[7296]  = 1;
  ram[7297]  = 1;
  ram[7298]  = 1;
  ram[7299]  = 1;
  ram[7300]  = 1;
  ram[7301]  = 1;
  ram[7302]  = 1;
  ram[7303]  = 1;
  ram[7304]  = 1;
  ram[7305]  = 1;
  ram[7306]  = 1;
  ram[7307]  = 1;
  ram[7308]  = 1;
  ram[7309]  = 1;
  ram[7310]  = 1;
  ram[7311]  = 1;
  ram[7312]  = 1;
  ram[7313]  = 1;
  ram[7314]  = 1;
  ram[7315]  = 0;
  ram[7316]  = 0;
  ram[7317]  = 0;
  ram[7318]  = 0;
  ram[7319]  = 0;
  ram[7320]  = 0;
  ram[7321]  = 0;
  ram[7322]  = 0;
  ram[7323]  = 0;
  ram[7324]  = 0;
  ram[7325]  = 0;
  ram[7326]  = 0;
  ram[7327]  = 1;
  ram[7328]  = 1;
  ram[7329]  = 1;
  ram[7330]  = 1;
  ram[7331]  = 0;
  ram[7332]  = 0;
  ram[7333]  = 0;
  ram[7334]  = 1;
  ram[7335]  = 1;
  ram[7336]  = 1;
  ram[7337]  = 1;
  ram[7338]  = 1;
  ram[7339]  = 1;
  ram[7340]  = 1;
  ram[7341]  = 1;
  ram[7342]  = 0;
  ram[7343]  = 0;
  ram[7344]  = 0;
  ram[7345]  = 1;
  ram[7346]  = 1;
  ram[7347]  = 1;
  ram[7348]  = 1;
  ram[7349]  = 1;
  ram[7350]  = 1;
  ram[7351]  = 1;
  ram[7352]  = 1;
  ram[7353]  = 1;
  ram[7354]  = 1;
  ram[7355]  = 1;
  ram[7356]  = 1;
  ram[7357]  = 1;
  ram[7358]  = 1;
  ram[7359]  = 1;
  ram[7360]  = 1;
  ram[7361]  = 1;
  ram[7362]  = 1;
  ram[7363]  = 1;
  ram[7364]  = 1;
  ram[7365]  = 1;
  ram[7366]  = 1;
  ram[7367]  = 1;
  ram[7368]  = 1;
  ram[7369]  = 1;
  ram[7370]  = 1;
  ram[7371]  = 1;
  ram[7372]  = 1;
  ram[7373]  = 1;
  ram[7374]  = 1;
  ram[7375]  = 1;
  ram[7376]  = 1;
  ram[7377]  = 1;
  ram[7378]  = 0;
  ram[7379]  = 0;
  ram[7380]  = 0;
  ram[7381]  = 0;
  ram[7382]  = 0;
  ram[7383]  = 1;
  ram[7384]  = 1;
  ram[7385]  = 1;
  ram[7386]  = 1;
  ram[7387]  = 1;
  ram[7388]  = 1;
  ram[7389]  = 1;
  ram[7390]  = 1;
  ram[7391]  = 1;
  ram[7392]  = 1;
  ram[7393]  = 1;
  ram[7394]  = 1;
  ram[7395]  = 1;
  ram[7396]  = 1;
  ram[7397]  = 1;
  ram[7398]  = 1;
  ram[7399]  = 1;
  ram[7400]  = 1;
  ram[7401]  = 1;
  ram[7402]  = 1;
  ram[7403]  = 1;
  ram[7404]  = 1;
  ram[7405]  = 1;
  ram[7406]  = 1;
  ram[7407]  = 1;
  ram[7408]  = 1;
  ram[7409]  = 1;
  ram[7410]  = 1;
  ram[7411]  = 1;
  ram[7412]  = 1;
  ram[7413]  = 1;
  ram[7414]  = 1;
  ram[7415]  = 1;
  ram[7416]  = 1;
  ram[7417]  = 1;
  ram[7418]  = 1;
  ram[7419]  = 1;
  ram[7420]  = 0;
  ram[7421]  = 0;
  ram[7422]  = 1;
  ram[7423]  = 1;
  ram[7424]  = 1;
  ram[7425]  = 1;
  ram[7426]  = 0;
  ram[7427]  = 0;
  ram[7428]  = 1;
  ram[7429]  = 1;
  ram[7430]  = 1;
  ram[7431]  = 1;
  ram[7432]  = 1;
  ram[7433]  = 1;
  ram[7434]  = 1;
  ram[7435]  = 0;
  ram[7436]  = 1;
  ram[7437]  = 1;
  ram[7438]  = 1;
  ram[7439]  = 1;
  ram[7440]  = 1;
  ram[7441]  = 1;
  ram[7442]  = 1;
  ram[7443]  = 0;
  ram[7444]  = 0;
  ram[7445]  = 1;
  ram[7446]  = 1;
  ram[7447]  = 1;
  ram[7448]  = 1;
  ram[7449]  = 1;
  ram[7450]  = 1;
  ram[7451]  = 1;
  ram[7452]  = 1;
  ram[7453]  = 1;
  ram[7454]  = 1;
  ram[7455]  = 1;
  ram[7456]  = 1;
  ram[7457]  = 0;
  ram[7458]  = 0;
  ram[7459]  = 1;
  ram[7460]  = 1;
  ram[7461]  = 1;
  ram[7462]  = 1;
  ram[7463]  = 1;
  ram[7464]  = 0;
  ram[7465]  = 0;
  ram[7466]  = 1;
  ram[7467]  = 1;
  ram[7468]  = 1;
  ram[7469]  = 1;
  ram[7470]  = 1;
  ram[7471]  = 1;
  ram[7472]  = 1;
  ram[7473]  = 1;
  ram[7474]  = 1;
  ram[7475]  = 0;
  ram[7476]  = 0;
  ram[7477]  = 1;
  ram[7478]  = 1;
  ram[7479]  = 1;
  ram[7480]  = 1;
  ram[7481]  = 0;
  ram[7482]  = 0;
  ram[7483]  = 1;
  ram[7484]  = 1;
  ram[7485]  = 1;
  ram[7486]  = 1;
  ram[7487]  = 1;
  ram[7488]  = 1;
  ram[7489]  = 1;
  ram[7490]  = 1;
  ram[7491]  = 1;
  ram[7492]  = 1;
  ram[7493]  = 1;
  ram[7494]  = 1;
  ram[7495]  = 1;
  ram[7496]  = 1;
  ram[7497]  = 1;
  ram[7498]  = 1;
  ram[7499]  = 1;
  ram[7500]  = 1;
  ram[7501]  = 1;
  ram[7502]  = 1;
  ram[7503]  = 1;
  ram[7504]  = 1;
  ram[7505]  = 1;
  ram[7506]  = 1;
  ram[7507]  = 1;
  ram[7508]  = 1;
  ram[7509]  = 1;
  ram[7510]  = 1;
  ram[7511]  = 1;
  ram[7512]  = 1;
  ram[7513]  = 1;
  ram[7514]  = 1;
  ram[7515]  = 1;
  ram[7516]  = 1;
  ram[7517]  = 1;
  ram[7518]  = 0;
  ram[7519]  = 0;
  ram[7520]  = 1;
  ram[7521]  = 1;
  ram[7522]  = 1;
  ram[7523]  = 1;
  ram[7524]  = 1;
  ram[7525]  = 1;
  ram[7526]  = 1;
  ram[7527]  = 1;
  ram[7528]  = 1;
  ram[7529]  = 1;
  ram[7530]  = 0;
  ram[7531]  = 0;
  ram[7532]  = 0;
  ram[7533]  = 1;
  ram[7534]  = 1;
  ram[7535]  = 1;
  ram[7536]  = 1;
  ram[7537]  = 1;
  ram[7538]  = 1;
  ram[7539]  = 1;
  ram[7540]  = 1;
  ram[7541]  = 1;
  ram[7542]  = 1;
  ram[7543]  = 0;
  ram[7544]  = 0;
  ram[7545]  = 0;
  ram[7546]  = 1;
  ram[7547]  = 1;
  ram[7548]  = 1;
  ram[7549]  = 1;
  ram[7550]  = 1;
  ram[7551]  = 1;
  ram[7552]  = 1;
  ram[7553]  = 1;
  ram[7554]  = 1;
  ram[7555]  = 1;
  ram[7556]  = 1;
  ram[7557]  = 1;
  ram[7558]  = 1;
  ram[7559]  = 1;
  ram[7560]  = 1;
  ram[7561]  = 1;
  ram[7562]  = 1;
  ram[7563]  = 1;
  ram[7564]  = 1;
  ram[7565]  = 1;
  ram[7566]  = 1;
  ram[7567]  = 1;
  ram[7568]  = 1;
  ram[7569]  = 1;
  ram[7570]  = 1;
  ram[7571]  = 1;
  ram[7572]  = 1;
  ram[7573]  = 1;
  ram[7574]  = 1;
  ram[7575]  = 1;
  ram[7576]  = 1;
  ram[7577]  = 0;
  ram[7578]  = 0;
  ram[7579]  = 0;
  ram[7580]  = 0;
  ram[7581]  = 1;
  ram[7582]  = 1;
  ram[7583]  = 1;
  ram[7584]  = 1;
  ram[7585]  = 1;
  ram[7586]  = 1;
  ram[7587]  = 1;
  ram[7588]  = 1;
  ram[7589]  = 1;
  ram[7590]  = 1;
  ram[7591]  = 1;
  ram[7592]  = 1;
  ram[7593]  = 1;
  ram[7594]  = 1;
  ram[7595]  = 1;
  ram[7596]  = 1;
  ram[7597]  = 1;
  ram[7598]  = 1;
  ram[7599]  = 1;
  ram[7600]  = 1;
  ram[7601]  = 1;
  ram[7602]  = 1;
  ram[7603]  = 1;
  ram[7604]  = 1;
  ram[7605]  = 1;
  ram[7606]  = 1;
  ram[7607]  = 1;
  ram[7608]  = 1;
  ram[7609]  = 1;
  ram[7610]  = 1;
  ram[7611]  = 1;
  ram[7612]  = 1;
  ram[7613]  = 1;
  ram[7614]  = 1;
  ram[7615]  = 1;
  ram[7616]  = 1;
  ram[7617]  = 1;
  ram[7618]  = 1;
  ram[7619]  = 1;
  ram[7620]  = 0;
  ram[7621]  = 0;
  ram[7622]  = 1;
  ram[7623]  = 1;
  ram[7624]  = 1;
  ram[7625]  = 1;
  ram[7626]  = 0;
  ram[7627]  = 0;
  ram[7628]  = 1;
  ram[7629]  = 1;
  ram[7630]  = 1;
  ram[7631]  = 1;
  ram[7632]  = 1;
  ram[7633]  = 1;
  ram[7634]  = 1;
  ram[7635]  = 0;
  ram[7636]  = 1;
  ram[7637]  = 1;
  ram[7638]  = 1;
  ram[7639]  = 1;
  ram[7640]  = 1;
  ram[7641]  = 1;
  ram[7642]  = 1;
  ram[7643]  = 0;
  ram[7644]  = 0;
  ram[7645]  = 1;
  ram[7646]  = 1;
  ram[7647]  = 1;
  ram[7648]  = 1;
  ram[7649]  = 1;
  ram[7650]  = 1;
  ram[7651]  = 1;
  ram[7652]  = 1;
  ram[7653]  = 1;
  ram[7654]  = 1;
  ram[7655]  = 1;
  ram[7656]  = 1;
  ram[7657]  = 0;
  ram[7658]  = 0;
  ram[7659]  = 1;
  ram[7660]  = 1;
  ram[7661]  = 1;
  ram[7662]  = 1;
  ram[7663]  = 1;
  ram[7664]  = 0;
  ram[7665]  = 0;
  ram[7666]  = 1;
  ram[7667]  = 1;
  ram[7668]  = 1;
  ram[7669]  = 1;
  ram[7670]  = 1;
  ram[7671]  = 1;
  ram[7672]  = 1;
  ram[7673]  = 1;
  ram[7674]  = 0;
  ram[7675]  = 0;
  ram[7676]  = 0;
  ram[7677]  = 1;
  ram[7678]  = 1;
  ram[7679]  = 1;
  ram[7680]  = 1;
  ram[7681]  = 0;
  ram[7682]  = 0;
  ram[7683]  = 1;
  ram[7684]  = 1;
  ram[7685]  = 1;
  ram[7686]  = 1;
  ram[7687]  = 1;
  ram[7688]  = 1;
  ram[7689]  = 1;
  ram[7690]  = 1;
  ram[7691]  = 1;
  ram[7692]  = 1;
  ram[7693]  = 1;
  ram[7694]  = 1;
  ram[7695]  = 1;
  ram[7696]  = 1;
  ram[7697]  = 1;
  ram[7698]  = 1;
  ram[7699]  = 1;
  ram[7700]  = 1;
  ram[7701]  = 1;
  ram[7702]  = 1;
  ram[7703]  = 1;
  ram[7704]  = 1;
  ram[7705]  = 1;
  ram[7706]  = 1;
  ram[7707]  = 1;
  ram[7708]  = 1;
  ram[7709]  = 1;
  ram[7710]  = 1;
  ram[7711]  = 1;
  ram[7712]  = 1;
  ram[7713]  = 1;
  ram[7714]  = 1;
  ram[7715]  = 1;
  ram[7716]  = 1;
  ram[7717]  = 1;
  ram[7718]  = 0;
  ram[7719]  = 1;
  ram[7720]  = 1;
  ram[7721]  = 1;
  ram[7722]  = 1;
  ram[7723]  = 1;
  ram[7724]  = 1;
  ram[7725]  = 1;
  ram[7726]  = 1;
  ram[7727]  = 1;
  ram[7728]  = 0;
  ram[7729]  = 0;
  ram[7730]  = 0;
  ram[7731]  = 0;
  ram[7732]  = 1;
  ram[7733]  = 1;
  ram[7734]  = 1;
  ram[7735]  = 1;
  ram[7736]  = 1;
  ram[7737]  = 1;
  ram[7738]  = 1;
  ram[7739]  = 1;
  ram[7740]  = 1;
  ram[7741]  = 1;
  ram[7742]  = 1;
  ram[7743]  = 0;
  ram[7744]  = 0;
  ram[7745]  = 0;
  ram[7746]  = 0;
  ram[7747]  = 1;
  ram[7748]  = 1;
  ram[7749]  = 1;
  ram[7750]  = 1;
  ram[7751]  = 1;
  ram[7752]  = 1;
  ram[7753]  = 1;
  ram[7754]  = 1;
  ram[7755]  = 1;
  ram[7756]  = 1;
  ram[7757]  = 1;
  ram[7758]  = 1;
  ram[7759]  = 1;
  ram[7760]  = 1;
  ram[7761]  = 1;
  ram[7762]  = 1;
  ram[7763]  = 1;
  ram[7764]  = 1;
  ram[7765]  = 1;
  ram[7766]  = 1;
  ram[7767]  = 1;
  ram[7768]  = 1;
  ram[7769]  = 1;
  ram[7770]  = 1;
  ram[7771]  = 1;
  ram[7772]  = 1;
  ram[7773]  = 1;
  ram[7774]  = 1;
  ram[7775]  = 0;
  ram[7776]  = 0;
  ram[7777]  = 0;
  ram[7778]  = 0;
  ram[7779]  = 0;
  ram[7780]  = 1;
  ram[7781]  = 1;
  ram[7782]  = 1;
  ram[7783]  = 1;
  ram[7784]  = 1;
  ram[7785]  = 1;
  ram[7786]  = 1;
  ram[7787]  = 1;
  ram[7788]  = 1;
  ram[7789]  = 1;
  ram[7790]  = 1;
  ram[7791]  = 1;
  ram[7792]  = 1;
  ram[7793]  = 1;
  ram[7794]  = 1;
  ram[7795]  = 1;
  ram[7796]  = 1;
  ram[7797]  = 1;
  ram[7798]  = 1;
  ram[7799]  = 1;
  ram[7800]  = 1;
  ram[7801]  = 1;
  ram[7802]  = 1;
  ram[7803]  = 1;
  ram[7804]  = 1;
  ram[7805]  = 1;
  ram[7806]  = 1;
  ram[7807]  = 1;
  ram[7808]  = 1;
  ram[7809]  = 1;
  ram[7810]  = 1;
  ram[7811]  = 1;
  ram[7812]  = 1;
  ram[7813]  = 1;
  ram[7814]  = 1;
  ram[7815]  = 1;
  ram[7816]  = 1;
  ram[7817]  = 1;
  ram[7818]  = 1;
  ram[7819]  = 1;
  ram[7820]  = 0;
  ram[7821]  = 0;
  ram[7822]  = 1;
  ram[7823]  = 1;
  ram[7824]  = 1;
  ram[7825]  = 1;
  ram[7826]  = 0;
  ram[7827]  = 0;
  ram[7828]  = 1;
  ram[7829]  = 1;
  ram[7830]  = 1;
  ram[7831]  = 1;
  ram[7832]  = 1;
  ram[7833]  = 1;
  ram[7834]  = 1;
  ram[7835]  = 0;
  ram[7836]  = 1;
  ram[7837]  = 1;
  ram[7838]  = 1;
  ram[7839]  = 1;
  ram[7840]  = 1;
  ram[7841]  = 1;
  ram[7842]  = 1;
  ram[7843]  = 0;
  ram[7844]  = 0;
  ram[7845]  = 1;
  ram[7846]  = 1;
  ram[7847]  = 1;
  ram[7848]  = 1;
  ram[7849]  = 1;
  ram[7850]  = 1;
  ram[7851]  = 1;
  ram[7852]  = 1;
  ram[7853]  = 1;
  ram[7854]  = 1;
  ram[7855]  = 1;
  ram[7856]  = 1;
  ram[7857]  = 0;
  ram[7858]  = 0;
  ram[7859]  = 1;
  ram[7860]  = 1;
  ram[7861]  = 1;
  ram[7862]  = 1;
  ram[7863]  = 1;
  ram[7864]  = 0;
  ram[7865]  = 0;
  ram[7866]  = 1;
  ram[7867]  = 1;
  ram[7868]  = 1;
  ram[7869]  = 1;
  ram[7870]  = 1;
  ram[7871]  = 1;
  ram[7872]  = 1;
  ram[7873]  = 1;
  ram[7874]  = 0;
  ram[7875]  = 0;
  ram[7876]  = 1;
  ram[7877]  = 1;
  ram[7878]  = 1;
  ram[7879]  = 1;
  ram[7880]  = 1;
  ram[7881]  = 0;
  ram[7882]  = 0;
  ram[7883]  = 1;
  ram[7884]  = 1;
  ram[7885]  = 1;
  ram[7886]  = 1;
  ram[7887]  = 1;
  ram[7888]  = 1;
  ram[7889]  = 1;
  ram[7890]  = 1;
  ram[7891]  = 1;
  ram[7892]  = 1;
  ram[7893]  = 1;
  ram[7894]  = 1;
  ram[7895]  = 1;
  ram[7896]  = 1;
  ram[7897]  = 1;
  ram[7898]  = 1;
  ram[7899]  = 1;
  ram[7900]  = 1;
  ram[7901]  = 1;
  ram[7902]  = 1;
  ram[7903]  = 1;
  ram[7904]  = 1;
  ram[7905]  = 1;
  ram[7906]  = 1;
  ram[7907]  = 1;
  ram[7908]  = 1;
  ram[7909]  = 1;
  ram[7910]  = 1;
  ram[7911]  = 1;
  ram[7912]  = 1;
  ram[7913]  = 1;
  ram[7914]  = 1;
  ram[7915]  = 1;
  ram[7916]  = 1;
  ram[7917]  = 0;
  ram[7918]  = 0;
  ram[7919]  = 1;
  ram[7920]  = 1;
  ram[7921]  = 1;
  ram[7922]  = 1;
  ram[7923]  = 1;
  ram[7924]  = 1;
  ram[7925]  = 1;
  ram[7926]  = 1;
  ram[7927]  = 0;
  ram[7928]  = 0;
  ram[7929]  = 0;
  ram[7930]  = 1;
  ram[7931]  = 1;
  ram[7932]  = 0;
  ram[7933]  = 0;
  ram[7934]  = 0;
  ram[7935]  = 0;
  ram[7936]  = 0;
  ram[7937]  = 0;
  ram[7938]  = 0;
  ram[7939]  = 0;
  ram[7940]  = 0;
  ram[7941]  = 0;
  ram[7942]  = 0;
  ram[7943]  = 0;
  ram[7944]  = 1;
  ram[7945]  = 0;
  ram[7946]  = 0;
  ram[7947]  = 0;
  ram[7948]  = 0;
  ram[7949]  = 1;
  ram[7950]  = 1;
  ram[7951]  = 1;
  ram[7952]  = 1;
  ram[7953]  = 1;
  ram[7954]  = 1;
  ram[7955]  = 1;
  ram[7956]  = 1;
  ram[7957]  = 1;
  ram[7958]  = 1;
  ram[7959]  = 1;
  ram[7960]  = 1;
  ram[7961]  = 1;
  ram[7962]  = 1;
  ram[7963]  = 1;
  ram[7964]  = 1;
  ram[7965]  = 1;
  ram[7966]  = 1;
  ram[7967]  = 1;
  ram[7968]  = 1;
  ram[7969]  = 1;
  ram[7970]  = 1;
  ram[7971]  = 1;
  ram[7972]  = 1;
  ram[7973]  = 1;
  ram[7974]  = 0;
  ram[7975]  = 0;
  ram[7976]  = 0;
  ram[7977]  = 0;
  ram[7978]  = 1;
  ram[7979]  = 1;
  ram[7980]  = 1;
  ram[7981]  = 1;
  ram[7982]  = 1;
  ram[7983]  = 1;
  ram[7984]  = 1;
  ram[7985]  = 1;
  ram[7986]  = 1;
  ram[7987]  = 1;
  ram[7988]  = 1;
  ram[7989]  = 1;
  ram[7990]  = 1;
  ram[7991]  = 1;
  ram[7992]  = 1;
  ram[7993]  = 1;
  ram[7994]  = 1;
  ram[7995]  = 1;
  ram[7996]  = 1;
  ram[7997]  = 1;
  ram[7998]  = 1;
  ram[7999]  = 1;
  ram[8000]  = 1;
  ram[8001]  = 1;
  ram[8002]  = 1;
  ram[8003]  = 1;
  ram[8004]  = 1;
  ram[8005]  = 1;
  ram[8006]  = 1;
  ram[8007]  = 1;
  ram[8008]  = 1;
  ram[8009]  = 1;
  ram[8010]  = 1;
  ram[8011]  = 1;
  ram[8012]  = 1;
  ram[8013]  = 1;
  ram[8014]  = 1;
  ram[8015]  = 1;
  ram[8016]  = 1;
  ram[8017]  = 1;
  ram[8018]  = 1;
  ram[8019]  = 1;
  ram[8020]  = 0;
  ram[8021]  = 0;
  ram[8022]  = 1;
  ram[8023]  = 1;
  ram[8024]  = 1;
  ram[8025]  = 1;
  ram[8026]  = 0;
  ram[8027]  = 0;
  ram[8028]  = 1;
  ram[8029]  = 1;
  ram[8030]  = 1;
  ram[8031]  = 1;
  ram[8032]  = 1;
  ram[8033]  = 1;
  ram[8034]  = 1;
  ram[8035]  = 0;
  ram[8036]  = 1;
  ram[8037]  = 1;
  ram[8038]  = 1;
  ram[8039]  = 1;
  ram[8040]  = 1;
  ram[8041]  = 1;
  ram[8042]  = 1;
  ram[8043]  = 0;
  ram[8044]  = 0;
  ram[8045]  = 1;
  ram[8046]  = 1;
  ram[8047]  = 1;
  ram[8048]  = 1;
  ram[8049]  = 1;
  ram[8050]  = 1;
  ram[8051]  = 1;
  ram[8052]  = 1;
  ram[8053]  = 1;
  ram[8054]  = 1;
  ram[8055]  = 1;
  ram[8056]  = 1;
  ram[8057]  = 0;
  ram[8058]  = 0;
  ram[8059]  = 1;
  ram[8060]  = 1;
  ram[8061]  = 1;
  ram[8062]  = 1;
  ram[8063]  = 1;
  ram[8064]  = 0;
  ram[8065]  = 0;
  ram[8066]  = 1;
  ram[8067]  = 1;
  ram[8068]  = 1;
  ram[8069]  = 1;
  ram[8070]  = 1;
  ram[8071]  = 1;
  ram[8072]  = 1;
  ram[8073]  = 0;
  ram[8074]  = 0;
  ram[8075]  = 1;
  ram[8076]  = 1;
  ram[8077]  = 1;
  ram[8078]  = 1;
  ram[8079]  = 1;
  ram[8080]  = 1;
  ram[8081]  = 0;
  ram[8082]  = 0;
  ram[8083]  = 1;
  ram[8084]  = 1;
  ram[8085]  = 1;
  ram[8086]  = 1;
  ram[8087]  = 1;
  ram[8088]  = 1;
  ram[8089]  = 1;
  ram[8090]  = 1;
  ram[8091]  = 1;
  ram[8092]  = 1;
  ram[8093]  = 1;
  ram[8094]  = 1;
  ram[8095]  = 1;
  ram[8096]  = 1;
  ram[8097]  = 1;
  ram[8098]  = 1;
  ram[8099]  = 1;
  ram[8100]  = 1;
  ram[8101]  = 1;
  ram[8102]  = 1;
  ram[8103]  = 1;
  ram[8104]  = 1;
  ram[8105]  = 1;
  ram[8106]  = 1;
  ram[8107]  = 1;
  ram[8108]  = 1;
  ram[8109]  = 1;
  ram[8110]  = 1;
  ram[8111]  = 1;
  ram[8112]  = 1;
  ram[8113]  = 1;
  ram[8114]  = 1;
  ram[8115]  = 1;
  ram[8116]  = 1;
  ram[8117]  = 0;
  ram[8118]  = 0;
  ram[8119]  = 1;
  ram[8120]  = 1;
  ram[8121]  = 1;
  ram[8122]  = 1;
  ram[8123]  = 1;
  ram[8124]  = 1;
  ram[8125]  = 1;
  ram[8126]  = 0;
  ram[8127]  = 0;
  ram[8128]  = 0;
  ram[8129]  = 1;
  ram[8130]  = 1;
  ram[8131]  = 1;
  ram[8132]  = 1;
  ram[8133]  = 1;
  ram[8134]  = 1;
  ram[8135]  = 1;
  ram[8136]  = 1;
  ram[8137]  = 1;
  ram[8138]  = 1;
  ram[8139]  = 1;
  ram[8140]  = 1;
  ram[8141]  = 1;
  ram[8142]  = 1;
  ram[8143]  = 1;
  ram[8144]  = 1;
  ram[8145]  = 1;
  ram[8146]  = 1;
  ram[8147]  = 0;
  ram[8148]  = 0;
  ram[8149]  = 1;
  ram[8150]  = 1;
  ram[8151]  = 1;
  ram[8152]  = 1;
  ram[8153]  = 1;
  ram[8154]  = 1;
  ram[8155]  = 1;
  ram[8156]  = 1;
  ram[8157]  = 1;
  ram[8158]  = 1;
  ram[8159]  = 1;
  ram[8160]  = 1;
  ram[8161]  = 1;
  ram[8162]  = 1;
  ram[8163]  = 1;
  ram[8164]  = 1;
  ram[8165]  = 1;
  ram[8166]  = 1;
  ram[8167]  = 1;
  ram[8168]  = 1;
  ram[8169]  = 1;
  ram[8170]  = 1;
  ram[8171]  = 1;
  ram[8172]  = 0;
  ram[8173]  = 0;
  ram[8174]  = 0;
  ram[8175]  = 0;
  ram[8176]  = 0;
  ram[8177]  = 1;
  ram[8178]  = 1;
  ram[8179]  = 1;
  ram[8180]  = 1;
  ram[8181]  = 1;
  ram[8182]  = 1;
  ram[8183]  = 1;
  ram[8184]  = 1;
  ram[8185]  = 1;
  ram[8186]  = 1;
  ram[8187]  = 1;
  ram[8188]  = 1;
  ram[8189]  = 1;
  ram[8190]  = 1;
  ram[8191]  = 1;
  ram[8192]  = 1;
  ram[8193]  = 1;
  ram[8194]  = 1;
  ram[8195]  = 1;
  ram[8196]  = 1;
  ram[8197]  = 1;
  ram[8198]  = 1;
  ram[8199]  = 1;
  ram[8200]  = 1;
  ram[8201]  = 1;
  ram[8202]  = 1;
  ram[8203]  = 1;
  ram[8204]  = 1;
  ram[8205]  = 1;
  ram[8206]  = 1;
  ram[8207]  = 1;
  ram[8208]  = 1;
  ram[8209]  = 1;
  ram[8210]  = 1;
  ram[8211]  = 1;
  ram[8212]  = 1;
  ram[8213]  = 1;
  ram[8214]  = 1;
  ram[8215]  = 1;
  ram[8216]  = 1;
  ram[8217]  = 1;
  ram[8218]  = 1;
  ram[8219]  = 1;
  ram[8220]  = 0;
  ram[8221]  = 0;
  ram[8222]  = 1;
  ram[8223]  = 1;
  ram[8224]  = 1;
  ram[8225]  = 1;
  ram[8226]  = 0;
  ram[8227]  = 0;
  ram[8228]  = 1;
  ram[8229]  = 0;
  ram[8230]  = 0;
  ram[8231]  = 0;
  ram[8232]  = 0;
  ram[8233]  = 0;
  ram[8234]  = 0;
  ram[8235]  = 0;
  ram[8236]  = 0;
  ram[8237]  = 0;
  ram[8238]  = 0;
  ram[8239]  = 0;
  ram[8240]  = 0;
  ram[8241]  = 0;
  ram[8242]  = 0;
  ram[8243]  = 0;
  ram[8244]  = 0;
  ram[8245]  = 0;
  ram[8246]  = 0;
  ram[8247]  = 0;
  ram[8248]  = 0;
  ram[8249]  = 0;
  ram[8250]  = 0;
  ram[8251]  = 0;
  ram[8252]  = 0;
  ram[8253]  = 1;
  ram[8254]  = 1;
  ram[8255]  = 1;
  ram[8256]  = 1;
  ram[8257]  = 0;
  ram[8258]  = 0;
  ram[8259]  = 1;
  ram[8260]  = 1;
  ram[8261]  = 1;
  ram[8262]  = 1;
  ram[8263]  = 1;
  ram[8264]  = 0;
  ram[8265]  = 0;
  ram[8266]  = 1;
  ram[8267]  = 1;
  ram[8268]  = 1;
  ram[8269]  = 1;
  ram[8270]  = 1;
  ram[8271]  = 1;
  ram[8272]  = 0;
  ram[8273]  = 0;
  ram[8274]  = 0;
  ram[8275]  = 1;
  ram[8276]  = 1;
  ram[8277]  = 1;
  ram[8278]  = 1;
  ram[8279]  = 1;
  ram[8280]  = 1;
  ram[8281]  = 0;
  ram[8282]  = 0;
  ram[8283]  = 1;
  ram[8284]  = 1;
  ram[8285]  = 1;
  ram[8286]  = 1;
  ram[8287]  = 1;
  ram[8288]  = 1;
  ram[8289]  = 1;
  ram[8290]  = 1;
  ram[8291]  = 1;
  ram[8292]  = 1;
  ram[8293]  = 1;
  ram[8294]  = 1;
  ram[8295]  = 1;
  ram[8296]  = 1;
  ram[8297]  = 1;
  ram[8298]  = 1;
  ram[8299]  = 1;
  ram[8300]  = 1;
  ram[8301]  = 1;
  ram[8302]  = 1;
  ram[8303]  = 1;
  ram[8304]  = 1;
  ram[8305]  = 1;
  ram[8306]  = 1;
  ram[8307]  = 1;
  ram[8308]  = 1;
  ram[8309]  = 1;
  ram[8310]  = 1;
  ram[8311]  = 1;
  ram[8312]  = 1;
  ram[8313]  = 1;
  ram[8314]  = 1;
  ram[8315]  = 1;
  ram[8316]  = 1;
  ram[8317]  = 0;
  ram[8318]  = 0;
  ram[8319]  = 1;
  ram[8320]  = 1;
  ram[8321]  = 0;
  ram[8322]  = 0;
  ram[8323]  = 1;
  ram[8324]  = 1;
  ram[8325]  = 1;
  ram[8326]  = 1;
  ram[8327]  = 0;
  ram[8328]  = 1;
  ram[8329]  = 1;
  ram[8330]  = 1;
  ram[8331]  = 1;
  ram[8332]  = 1;
  ram[8333]  = 1;
  ram[8334]  = 1;
  ram[8335]  = 1;
  ram[8336]  = 1;
  ram[8337]  = 1;
  ram[8338]  = 1;
  ram[8339]  = 1;
  ram[8340]  = 1;
  ram[8341]  = 1;
  ram[8342]  = 1;
  ram[8343]  = 1;
  ram[8344]  = 1;
  ram[8345]  = 1;
  ram[8346]  = 1;
  ram[8347]  = 1;
  ram[8348]  = 1;
  ram[8349]  = 1;
  ram[8350]  = 1;
  ram[8351]  = 1;
  ram[8352]  = 1;
  ram[8353]  = 1;
  ram[8354]  = 1;
  ram[8355]  = 1;
  ram[8356]  = 1;
  ram[8357]  = 1;
  ram[8358]  = 1;
  ram[8359]  = 1;
  ram[8360]  = 1;
  ram[8361]  = 1;
  ram[8362]  = 1;
  ram[8363]  = 1;
  ram[8364]  = 1;
  ram[8365]  = 1;
  ram[8366]  = 1;
  ram[8367]  = 1;
  ram[8368]  = 1;
  ram[8369]  = 1;
  ram[8370]  = 1;
  ram[8371]  = 0;
  ram[8372]  = 0;
  ram[8373]  = 0;
  ram[8374]  = 0;
  ram[8375]  = 1;
  ram[8376]  = 1;
  ram[8377]  = 1;
  ram[8378]  = 1;
  ram[8379]  = 1;
  ram[8380]  = 1;
  ram[8381]  = 1;
  ram[8382]  = 1;
  ram[8383]  = 1;
  ram[8384]  = 1;
  ram[8385]  = 1;
  ram[8386]  = 1;
  ram[8387]  = 1;
  ram[8388]  = 1;
  ram[8389]  = 1;
  ram[8390]  = 1;
  ram[8391]  = 1;
  ram[8392]  = 1;
  ram[8393]  = 1;
  ram[8394]  = 1;
  ram[8395]  = 1;
  ram[8396]  = 1;
  ram[8397]  = 1;
  ram[8398]  = 1;
  ram[8399]  = 1;
  ram[8400]  = 1;
  ram[8401]  = 1;
  ram[8402]  = 1;
  ram[8403]  = 1;
  ram[8404]  = 1;
  ram[8405]  = 1;
  ram[8406]  = 1;
  ram[8407]  = 1;
  ram[8408]  = 1;
  ram[8409]  = 1;
  ram[8410]  = 1;
  ram[8411]  = 1;
  ram[8412]  = 1;
  ram[8413]  = 1;
  ram[8414]  = 1;
  ram[8415]  = 1;
  ram[8416]  = 1;
  ram[8417]  = 1;
  ram[8418]  = 1;
  ram[8419]  = 1;
  ram[8420]  = 0;
  ram[8421]  = 0;
  ram[8422]  = 1;
  ram[8423]  = 1;
  ram[8424]  = 1;
  ram[8425]  = 1;
  ram[8426]  = 0;
  ram[8427]  = 0;
  ram[8428]  = 1;
  ram[8429]  = 0;
  ram[8430]  = 0;
  ram[8431]  = 0;
  ram[8432]  = 0;
  ram[8433]  = 0;
  ram[8434]  = 0;
  ram[8435]  = 0;
  ram[8436]  = 0;
  ram[8437]  = 0;
  ram[8438]  = 0;
  ram[8439]  = 0;
  ram[8440]  = 0;
  ram[8441]  = 0;
  ram[8442]  = 0;
  ram[8443]  = 0;
  ram[8444]  = 0;
  ram[8445]  = 0;
  ram[8446]  = 0;
  ram[8447]  = 0;
  ram[8448]  = 0;
  ram[8449]  = 0;
  ram[8450]  = 0;
  ram[8451]  = 0;
  ram[8452]  = 0;
  ram[8453]  = 1;
  ram[8454]  = 1;
  ram[8455]  = 1;
  ram[8456]  = 1;
  ram[8457]  = 0;
  ram[8458]  = 0;
  ram[8459]  = 1;
  ram[8460]  = 1;
  ram[8461]  = 1;
  ram[8462]  = 1;
  ram[8463]  = 1;
  ram[8464]  = 0;
  ram[8465]  = 0;
  ram[8466]  = 1;
  ram[8467]  = 1;
  ram[8468]  = 1;
  ram[8469]  = 1;
  ram[8470]  = 1;
  ram[8471]  = 1;
  ram[8472]  = 0;
  ram[8473]  = 0;
  ram[8474]  = 1;
  ram[8475]  = 1;
  ram[8476]  = 1;
  ram[8477]  = 1;
  ram[8478]  = 1;
  ram[8479]  = 1;
  ram[8480]  = 1;
  ram[8481]  = 0;
  ram[8482]  = 0;
  ram[8483]  = 1;
  ram[8484]  = 1;
  ram[8485]  = 1;
  ram[8486]  = 1;
  ram[8487]  = 1;
  ram[8488]  = 1;
  ram[8489]  = 1;
  ram[8490]  = 1;
  ram[8491]  = 1;
  ram[8492]  = 1;
  ram[8493]  = 1;
  ram[8494]  = 1;
  ram[8495]  = 1;
  ram[8496]  = 1;
  ram[8497]  = 1;
  ram[8498]  = 1;
  ram[8499]  = 1;
  ram[8500]  = 1;
  ram[8501]  = 1;
  ram[8502]  = 1;
  ram[8503]  = 1;
  ram[8504]  = 1;
  ram[8505]  = 1;
  ram[8506]  = 1;
  ram[8507]  = 1;
  ram[8508]  = 1;
  ram[8509]  = 1;
  ram[8510]  = 1;
  ram[8511]  = 1;
  ram[8512]  = 1;
  ram[8513]  = 1;
  ram[8514]  = 1;
  ram[8515]  = 1;
  ram[8516]  = 1;
  ram[8517]  = 0;
  ram[8518]  = 1;
  ram[8519]  = 1;
  ram[8520]  = 1;
  ram[8521]  = 0;
  ram[8522]  = 0;
  ram[8523]  = 1;
  ram[8524]  = 1;
  ram[8525]  = 1;
  ram[8526]  = 1;
  ram[8527]  = 1;
  ram[8528]  = 1;
  ram[8529]  = 1;
  ram[8530]  = 1;
  ram[8531]  = 1;
  ram[8532]  = 1;
  ram[8533]  = 1;
  ram[8534]  = 1;
  ram[8535]  = 1;
  ram[8536]  = 1;
  ram[8537]  = 1;
  ram[8538]  = 1;
  ram[8539]  = 1;
  ram[8540]  = 1;
  ram[8541]  = 1;
  ram[8542]  = 1;
  ram[8543]  = 1;
  ram[8544]  = 1;
  ram[8545]  = 1;
  ram[8546]  = 1;
  ram[8547]  = 1;
  ram[8548]  = 1;
  ram[8549]  = 1;
  ram[8550]  = 1;
  ram[8551]  = 1;
  ram[8552]  = 1;
  ram[8553]  = 1;
  ram[8554]  = 1;
  ram[8555]  = 1;
  ram[8556]  = 1;
  ram[8557]  = 1;
  ram[8558]  = 1;
  ram[8559]  = 1;
  ram[8560]  = 1;
  ram[8561]  = 1;
  ram[8562]  = 1;
  ram[8563]  = 1;
  ram[8564]  = 1;
  ram[8565]  = 1;
  ram[8566]  = 1;
  ram[8567]  = 1;
  ram[8568]  = 1;
  ram[8569]  = 0;
  ram[8570]  = 0;
  ram[8571]  = 0;
  ram[8572]  = 0;
  ram[8573]  = 1;
  ram[8574]  = 1;
  ram[8575]  = 1;
  ram[8576]  = 1;
  ram[8577]  = 1;
  ram[8578]  = 1;
  ram[8579]  = 1;
  ram[8580]  = 1;
  ram[8581]  = 1;
  ram[8582]  = 1;
  ram[8583]  = 1;
  ram[8584]  = 1;
  ram[8585]  = 1;
  ram[8586]  = 1;
  ram[8587]  = 1;
  ram[8588]  = 1;
  ram[8589]  = 1;
  ram[8590]  = 1;
  ram[8591]  = 1;
  ram[8592]  = 1;
  ram[8593]  = 1;
  ram[8594]  = 1;
  ram[8595]  = 1;
  ram[8596]  = 1;
  ram[8597]  = 1;
  ram[8598]  = 1;
  ram[8599]  = 1;
  ram[8600]  = 1;
  ram[8601]  = 1;
  ram[8602]  = 1;
  ram[8603]  = 1;
  ram[8604]  = 1;
  ram[8605]  = 1;
  ram[8606]  = 1;
  ram[8607]  = 1;
  ram[8608]  = 1;
  ram[8609]  = 1;
  ram[8610]  = 1;
  ram[8611]  = 1;
  ram[8612]  = 1;
  ram[8613]  = 1;
  ram[8614]  = 1;
  ram[8615]  = 1;
  ram[8616]  = 1;
  ram[8617]  = 1;
  ram[8618]  = 1;
  ram[8619]  = 1;
  ram[8620]  = 0;
  ram[8621]  = 0;
  ram[8622]  = 1;
  ram[8623]  = 1;
  ram[8624]  = 1;
  ram[8625]  = 1;
  ram[8626]  = 0;
  ram[8627]  = 0;
  ram[8628]  = 1;
  ram[8629]  = 1;
  ram[8630]  = 1;
  ram[8631]  = 1;
  ram[8632]  = 1;
  ram[8633]  = 1;
  ram[8634]  = 1;
  ram[8635]  = 0;
  ram[8636]  = 1;
  ram[8637]  = 1;
  ram[8638]  = 1;
  ram[8639]  = 1;
  ram[8640]  = 1;
  ram[8641]  = 1;
  ram[8642]  = 1;
  ram[8643]  = 0;
  ram[8644]  = 0;
  ram[8645]  = 1;
  ram[8646]  = 1;
  ram[8647]  = 1;
  ram[8648]  = 1;
  ram[8649]  = 1;
  ram[8650]  = 1;
  ram[8651]  = 1;
  ram[8652]  = 1;
  ram[8653]  = 1;
  ram[8654]  = 1;
  ram[8655]  = 1;
  ram[8656]  = 1;
  ram[8657]  = 0;
  ram[8658]  = 0;
  ram[8659]  = 1;
  ram[8660]  = 1;
  ram[8661]  = 1;
  ram[8662]  = 1;
  ram[8663]  = 1;
  ram[8664]  = 0;
  ram[8665]  = 0;
  ram[8666]  = 1;
  ram[8667]  = 1;
  ram[8668]  = 1;
  ram[8669]  = 1;
  ram[8670]  = 1;
  ram[8671]  = 1;
  ram[8672]  = 0;
  ram[8673]  = 0;
  ram[8674]  = 1;
  ram[8675]  = 1;
  ram[8676]  = 1;
  ram[8677]  = 1;
  ram[8678]  = 1;
  ram[8679]  = 1;
  ram[8680]  = 1;
  ram[8681]  = 0;
  ram[8682]  = 0;
  ram[8683]  = 1;
  ram[8684]  = 1;
  ram[8685]  = 1;
  ram[8686]  = 1;
  ram[8687]  = 1;
  ram[8688]  = 1;
  ram[8689]  = 1;
  ram[8690]  = 1;
  ram[8691]  = 1;
  ram[8692]  = 1;
  ram[8693]  = 1;
  ram[8694]  = 1;
  ram[8695]  = 1;
  ram[8696]  = 1;
  ram[8697]  = 1;
  ram[8698]  = 1;
  ram[8699]  = 1;
  ram[8700]  = 1;
  ram[8701]  = 1;
  ram[8702]  = 1;
  ram[8703]  = 1;
  ram[8704]  = 1;
  ram[8705]  = 1;
  ram[8706]  = 1;
  ram[8707]  = 1;
  ram[8708]  = 1;
  ram[8709]  = 1;
  ram[8710]  = 1;
  ram[8711]  = 1;
  ram[8712]  = 1;
  ram[8713]  = 1;
  ram[8714]  = 1;
  ram[8715]  = 1;
  ram[8716]  = 0;
  ram[8717]  = 0;
  ram[8718]  = 1;
  ram[8719]  = 1;
  ram[8720]  = 1;
  ram[8721]  = 0;
  ram[8722]  = 0;
  ram[8723]  = 1;
  ram[8724]  = 1;
  ram[8725]  = 1;
  ram[8726]  = 1;
  ram[8727]  = 1;
  ram[8728]  = 1;
  ram[8729]  = 1;
  ram[8730]  = 1;
  ram[8731]  = 1;
  ram[8732]  = 1;
  ram[8733]  = 1;
  ram[8734]  = 1;
  ram[8735]  = 1;
  ram[8736]  = 1;
  ram[8737]  = 1;
  ram[8738]  = 1;
  ram[8739]  = 1;
  ram[8740]  = 1;
  ram[8741]  = 1;
  ram[8742]  = 1;
  ram[8743]  = 1;
  ram[8744]  = 1;
  ram[8745]  = 1;
  ram[8746]  = 0;
  ram[8747]  = 0;
  ram[8748]  = 1;
  ram[8749]  = 1;
  ram[8750]  = 1;
  ram[8751]  = 1;
  ram[8752]  = 1;
  ram[8753]  = 1;
  ram[8754]  = 1;
  ram[8755]  = 1;
  ram[8756]  = 1;
  ram[8757]  = 1;
  ram[8758]  = 1;
  ram[8759]  = 1;
  ram[8760]  = 1;
  ram[8761]  = 1;
  ram[8762]  = 1;
  ram[8763]  = 1;
  ram[8764]  = 1;
  ram[8765]  = 1;
  ram[8766]  = 1;
  ram[8767]  = 1;
  ram[8768]  = 1;
  ram[8769]  = 0;
  ram[8770]  = 0;
  ram[8771]  = 0;
  ram[8772]  = 1;
  ram[8773]  = 1;
  ram[8774]  = 1;
  ram[8775]  = 1;
  ram[8776]  = 1;
  ram[8777]  = 1;
  ram[8778]  = 1;
  ram[8779]  = 1;
  ram[8780]  = 1;
  ram[8781]  = 1;
  ram[8782]  = 1;
  ram[8783]  = 1;
  ram[8784]  = 1;
  ram[8785]  = 1;
  ram[8786]  = 1;
  ram[8787]  = 1;
  ram[8788]  = 1;
  ram[8789]  = 1;
  ram[8790]  = 1;
  ram[8791]  = 1;
  ram[8792]  = 1;
  ram[8793]  = 1;
  ram[8794]  = 1;
  ram[8795]  = 1;
  ram[8796]  = 1;
  ram[8797]  = 1;
  ram[8798]  = 1;
  ram[8799]  = 1;
  ram[8800]  = 1;
  ram[8801]  = 1;
  ram[8802]  = 1;
  ram[8803]  = 1;
  ram[8804]  = 1;
  ram[8805]  = 1;
  ram[8806]  = 1;
  ram[8807]  = 1;
  ram[8808]  = 1;
  ram[8809]  = 1;
  ram[8810]  = 1;
  ram[8811]  = 1;
  ram[8812]  = 1;
  ram[8813]  = 1;
  ram[8814]  = 1;
  ram[8815]  = 1;
  ram[8816]  = 1;
  ram[8817]  = 1;
  ram[8818]  = 1;
  ram[8819]  = 1;
  ram[8820]  = 0;
  ram[8821]  = 0;
  ram[8822]  = 1;
  ram[8823]  = 1;
  ram[8824]  = 1;
  ram[8825]  = 1;
  ram[8826]  = 0;
  ram[8827]  = 0;
  ram[8828]  = 1;
  ram[8829]  = 1;
  ram[8830]  = 1;
  ram[8831]  = 1;
  ram[8832]  = 1;
  ram[8833]  = 1;
  ram[8834]  = 1;
  ram[8835]  = 0;
  ram[8836]  = 1;
  ram[8837]  = 1;
  ram[8838]  = 1;
  ram[8839]  = 1;
  ram[8840]  = 1;
  ram[8841]  = 1;
  ram[8842]  = 1;
  ram[8843]  = 0;
  ram[8844]  = 0;
  ram[8845]  = 1;
  ram[8846]  = 1;
  ram[8847]  = 1;
  ram[8848]  = 1;
  ram[8849]  = 1;
  ram[8850]  = 1;
  ram[8851]  = 1;
  ram[8852]  = 1;
  ram[8853]  = 1;
  ram[8854]  = 1;
  ram[8855]  = 1;
  ram[8856]  = 1;
  ram[8857]  = 0;
  ram[8858]  = 0;
  ram[8859]  = 1;
  ram[8860]  = 1;
  ram[8861]  = 1;
  ram[8862]  = 1;
  ram[8863]  = 1;
  ram[8864]  = 0;
  ram[8865]  = 0;
  ram[8866]  = 1;
  ram[8867]  = 1;
  ram[8868]  = 1;
  ram[8869]  = 1;
  ram[8870]  = 1;
  ram[8871]  = 1;
  ram[8872]  = 0;
  ram[8873]  = 0;
  ram[8874]  = 1;
  ram[8875]  = 1;
  ram[8876]  = 1;
  ram[8877]  = 1;
  ram[8878]  = 1;
  ram[8879]  = 1;
  ram[8880]  = 1;
  ram[8881]  = 0;
  ram[8882]  = 0;
  ram[8883]  = 1;
  ram[8884]  = 1;
  ram[8885]  = 1;
  ram[8886]  = 1;
  ram[8887]  = 1;
  ram[8888]  = 1;
  ram[8889]  = 1;
  ram[8890]  = 1;
  ram[8891]  = 1;
  ram[8892]  = 1;
  ram[8893]  = 1;
  ram[8894]  = 1;
  ram[8895]  = 1;
  ram[8896]  = 1;
  ram[8897]  = 1;
  ram[8898]  = 1;
  ram[8899]  = 1;
  ram[8900]  = 1;
  ram[8901]  = 1;
  ram[8902]  = 1;
  ram[8903]  = 1;
  ram[8904]  = 1;
  ram[8905]  = 1;
  ram[8906]  = 1;
  ram[8907]  = 1;
  ram[8908]  = 1;
  ram[8909]  = 1;
  ram[8910]  = 1;
  ram[8911]  = 1;
  ram[8912]  = 1;
  ram[8913]  = 1;
  ram[8914]  = 1;
  ram[8915]  = 1;
  ram[8916]  = 0;
  ram[8917]  = 0;
  ram[8918]  = 1;
  ram[8919]  = 1;
  ram[8920]  = 1;
  ram[8921]  = 0;
  ram[8922]  = 0;
  ram[8923]  = 1;
  ram[8924]  = 1;
  ram[8925]  = 1;
  ram[8926]  = 1;
  ram[8927]  = 1;
  ram[8928]  = 0;
  ram[8929]  = 0;
  ram[8930]  = 0;
  ram[8931]  = 0;
  ram[8932]  = 0;
  ram[8933]  = 0;
  ram[8934]  = 0;
  ram[8935]  = 0;
  ram[8936]  = 0;
  ram[8937]  = 1;
  ram[8938]  = 1;
  ram[8939]  = 1;
  ram[8940]  = 1;
  ram[8941]  = 1;
  ram[8942]  = 1;
  ram[8943]  = 1;
  ram[8944]  = 1;
  ram[8945]  = 1;
  ram[8946]  = 0;
  ram[8947]  = 0;
  ram[8948]  = 1;
  ram[8949]  = 1;
  ram[8950]  = 1;
  ram[8951]  = 1;
  ram[8952]  = 1;
  ram[8953]  = 1;
  ram[8954]  = 1;
  ram[8955]  = 1;
  ram[8956]  = 1;
  ram[8957]  = 1;
  ram[8958]  = 1;
  ram[8959]  = 1;
  ram[8960]  = 1;
  ram[8961]  = 1;
  ram[8962]  = 1;
  ram[8963]  = 1;
  ram[8964]  = 1;
  ram[8965]  = 1;
  ram[8966]  = 1;
  ram[8967]  = 1;
  ram[8968]  = 1;
  ram[8969]  = 0;
  ram[8970]  = 0;
  ram[8971]  = 1;
  ram[8972]  = 1;
  ram[8973]  = 1;
  ram[8974]  = 1;
  ram[8975]  = 1;
  ram[8976]  = 1;
  ram[8977]  = 1;
  ram[8978]  = 1;
  ram[8979]  = 1;
  ram[8980]  = 1;
  ram[8981]  = 1;
  ram[8982]  = 1;
  ram[8983]  = 1;
  ram[8984]  = 1;
  ram[8985]  = 1;
  ram[8986]  = 1;
  ram[8987]  = 1;
  ram[8988]  = 1;
  ram[8989]  = 1;
  ram[8990]  = 1;
  ram[8991]  = 1;
  ram[8992]  = 1;
  ram[8993]  = 1;
  ram[8994]  = 1;
  ram[8995]  = 1;
  ram[8996]  = 1;
  ram[8997]  = 1;
  ram[8998]  = 1;
  ram[8999]  = 1;
  ram[9000]  = 1;
  ram[9001]  = 1;
  ram[9002]  = 1;
  ram[9003]  = 1;
  ram[9004]  = 1;
  ram[9005]  = 1;
  ram[9006]  = 1;
  ram[9007]  = 1;
  ram[9008]  = 1;
  ram[9009]  = 1;
  ram[9010]  = 1;
  ram[9011]  = 1;
  ram[9012]  = 1;
  ram[9013]  = 1;
  ram[9014]  = 1;
  ram[9015]  = 1;
  ram[9016]  = 1;
  ram[9017]  = 1;
  ram[9018]  = 1;
  ram[9019]  = 1;
  ram[9020]  = 0;
  ram[9021]  = 0;
  ram[9022]  = 1;
  ram[9023]  = 1;
  ram[9024]  = 1;
  ram[9025]  = 1;
  ram[9026]  = 0;
  ram[9027]  = 0;
  ram[9028]  = 1;
  ram[9029]  = 1;
  ram[9030]  = 1;
  ram[9031]  = 1;
  ram[9032]  = 1;
  ram[9033]  = 1;
  ram[9034]  = 1;
  ram[9035]  = 0;
  ram[9036]  = 1;
  ram[9037]  = 1;
  ram[9038]  = 1;
  ram[9039]  = 1;
  ram[9040]  = 1;
  ram[9041]  = 1;
  ram[9042]  = 1;
  ram[9043]  = 0;
  ram[9044]  = 0;
  ram[9045]  = 1;
  ram[9046]  = 1;
  ram[9047]  = 1;
  ram[9048]  = 1;
  ram[9049]  = 1;
  ram[9050]  = 1;
  ram[9051]  = 1;
  ram[9052]  = 1;
  ram[9053]  = 1;
  ram[9054]  = 1;
  ram[9055]  = 1;
  ram[9056]  = 1;
  ram[9057]  = 0;
  ram[9058]  = 0;
  ram[9059]  = 1;
  ram[9060]  = 1;
  ram[9061]  = 1;
  ram[9062]  = 1;
  ram[9063]  = 1;
  ram[9064]  = 0;
  ram[9065]  = 0;
  ram[9066]  = 1;
  ram[9067]  = 1;
  ram[9068]  = 1;
  ram[9069]  = 1;
  ram[9070]  = 1;
  ram[9071]  = 1;
  ram[9072]  = 0;
  ram[9073]  = 0;
  ram[9074]  = 0;
  ram[9075]  = 0;
  ram[9076]  = 0;
  ram[9077]  = 0;
  ram[9078]  = 1;
  ram[9079]  = 1;
  ram[9080]  = 1;
  ram[9081]  = 0;
  ram[9082]  = 0;
  ram[9083]  = 1;
  ram[9084]  = 1;
  ram[9085]  = 1;
  ram[9086]  = 1;
  ram[9087]  = 1;
  ram[9088]  = 1;
  ram[9089]  = 1;
  ram[9090]  = 1;
  ram[9091]  = 1;
  ram[9092]  = 1;
  ram[9093]  = 1;
  ram[9094]  = 1;
  ram[9095]  = 1;
  ram[9096]  = 1;
  ram[9097]  = 1;
  ram[9098]  = 1;
  ram[9099]  = 1;
  ram[9100]  = 1;
  ram[9101]  = 1;
  ram[9102]  = 1;
  ram[9103]  = 1;
  ram[9104]  = 1;
  ram[9105]  = 1;
  ram[9106]  = 1;
  ram[9107]  = 1;
  ram[9108]  = 1;
  ram[9109]  = 1;
  ram[9110]  = 1;
  ram[9111]  = 1;
  ram[9112]  = 1;
  ram[9113]  = 1;
  ram[9114]  = 1;
  ram[9115]  = 1;
  ram[9116]  = 0;
  ram[9117]  = 1;
  ram[9118]  = 1;
  ram[9119]  = 1;
  ram[9120]  = 1;
  ram[9121]  = 0;
  ram[9122]  = 0;
  ram[9123]  = 1;
  ram[9124]  = 1;
  ram[9125]  = 1;
  ram[9126]  = 1;
  ram[9127]  = 1;
  ram[9128]  = 0;
  ram[9129]  = 0;
  ram[9130]  = 1;
  ram[9131]  = 1;
  ram[9132]  = 1;
  ram[9133]  = 1;
  ram[9134]  = 1;
  ram[9135]  = 0;
  ram[9136]  = 0;
  ram[9137]  = 1;
  ram[9138]  = 1;
  ram[9139]  = 1;
  ram[9140]  = 1;
  ram[9141]  = 0;
  ram[9142]  = 1;
  ram[9143]  = 1;
  ram[9144]  = 1;
  ram[9145]  = 1;
  ram[9146]  = 0;
  ram[9147]  = 0;
  ram[9148]  = 1;
  ram[9149]  = 1;
  ram[9150]  = 1;
  ram[9151]  = 1;
  ram[9152]  = 1;
  ram[9153]  = 1;
  ram[9154]  = 1;
  ram[9155]  = 1;
  ram[9156]  = 1;
  ram[9157]  = 1;
  ram[9158]  = 1;
  ram[9159]  = 1;
  ram[9160]  = 1;
  ram[9161]  = 1;
  ram[9162]  = 1;
  ram[9163]  = 1;
  ram[9164]  = 1;
  ram[9165]  = 1;
  ram[9166]  = 1;
  ram[9167]  = 1;
  ram[9168]  = 1;
  ram[9169]  = 0;
  ram[9170]  = 0;
  ram[9171]  = 1;
  ram[9172]  = 1;
  ram[9173]  = 1;
  ram[9174]  = 1;
  ram[9175]  = 1;
  ram[9176]  = 1;
  ram[9177]  = 1;
  ram[9178]  = 1;
  ram[9179]  = 1;
  ram[9180]  = 1;
  ram[9181]  = 1;
  ram[9182]  = 1;
  ram[9183]  = 1;
  ram[9184]  = 1;
  ram[9185]  = 1;
  ram[9186]  = 1;
  ram[9187]  = 1;
  ram[9188]  = 1;
  ram[9189]  = 1;
  ram[9190]  = 1;
  ram[9191]  = 1;
  ram[9192]  = 1;
  ram[9193]  = 1;
  ram[9194]  = 1;
  ram[9195]  = 1;
  ram[9196]  = 1;
  ram[9197]  = 1;
  ram[9198]  = 1;
  ram[9199]  = 1;
  ram[9200]  = 1;
  ram[9201]  = 1;
  ram[9202]  = 1;
  ram[9203]  = 1;
  ram[9204]  = 1;
  ram[9205]  = 1;
  ram[9206]  = 1;
  ram[9207]  = 1;
  ram[9208]  = 1;
  ram[9209]  = 1;
  ram[9210]  = 1;
  ram[9211]  = 1;
  ram[9212]  = 1;
  ram[9213]  = 1;
  ram[9214]  = 1;
  ram[9215]  = 1;
  ram[9216]  = 1;
  ram[9217]  = 1;
  ram[9218]  = 1;
  ram[9219]  = 1;
  ram[9220]  = 0;
  ram[9221]  = 0;
  ram[9222]  = 1;
  ram[9223]  = 1;
  ram[9224]  = 1;
  ram[9225]  = 1;
  ram[9226]  = 0;
  ram[9227]  = 0;
  ram[9228]  = 1;
  ram[9229]  = 1;
  ram[9230]  = 1;
  ram[9231]  = 1;
  ram[9232]  = 1;
  ram[9233]  = 1;
  ram[9234]  = 1;
  ram[9235]  = 0;
  ram[9236]  = 1;
  ram[9237]  = 1;
  ram[9238]  = 1;
  ram[9239]  = 1;
  ram[9240]  = 1;
  ram[9241]  = 1;
  ram[9242]  = 1;
  ram[9243]  = 0;
  ram[9244]  = 0;
  ram[9245]  = 1;
  ram[9246]  = 1;
  ram[9247]  = 1;
  ram[9248]  = 1;
  ram[9249]  = 1;
  ram[9250]  = 1;
  ram[9251]  = 0;
  ram[9252]  = 1;
  ram[9253]  = 1;
  ram[9254]  = 1;
  ram[9255]  = 1;
  ram[9256]  = 1;
  ram[9257]  = 0;
  ram[9258]  = 0;
  ram[9259]  = 1;
  ram[9260]  = 1;
  ram[9261]  = 1;
  ram[9262]  = 1;
  ram[9263]  = 1;
  ram[9264]  = 0;
  ram[9265]  = 0;
  ram[9266]  = 1;
  ram[9267]  = 1;
  ram[9268]  = 1;
  ram[9269]  = 1;
  ram[9270]  = 1;
  ram[9271]  = 1;
  ram[9272]  = 0;
  ram[9273]  = 0;
  ram[9274]  = 0;
  ram[9275]  = 0;
  ram[9276]  = 0;
  ram[9277]  = 0;
  ram[9278]  = 1;
  ram[9279]  = 1;
  ram[9280]  = 1;
  ram[9281]  = 0;
  ram[9282]  = 0;
  ram[9283]  = 1;
  ram[9284]  = 1;
  ram[9285]  = 1;
  ram[9286]  = 1;
  ram[9287]  = 1;
  ram[9288]  = 1;
  ram[9289]  = 1;
  ram[9290]  = 1;
  ram[9291]  = 1;
  ram[9292]  = 1;
  ram[9293]  = 1;
  ram[9294]  = 1;
  ram[9295]  = 1;
  ram[9296]  = 1;
  ram[9297]  = 1;
  ram[9298]  = 1;
  ram[9299]  = 1;
  ram[9300]  = 1;
  ram[9301]  = 1;
  ram[9302]  = 1;
  ram[9303]  = 1;
  ram[9304]  = 1;
  ram[9305]  = 1;
  ram[9306]  = 1;
  ram[9307]  = 1;
  ram[9308]  = 1;
  ram[9309]  = 1;
  ram[9310]  = 1;
  ram[9311]  = 1;
  ram[9312]  = 1;
  ram[9313]  = 1;
  ram[9314]  = 1;
  ram[9315]  = 0;
  ram[9316]  = 0;
  ram[9317]  = 1;
  ram[9318]  = 1;
  ram[9319]  = 1;
  ram[9320]  = 1;
  ram[9321]  = 0;
  ram[9322]  = 0;
  ram[9323]  = 1;
  ram[9324]  = 1;
  ram[9325]  = 1;
  ram[9326]  = 1;
  ram[9327]  = 1;
  ram[9328]  = 0;
  ram[9329]  = 0;
  ram[9330]  = 1;
  ram[9331]  = 1;
  ram[9332]  = 1;
  ram[9333]  = 1;
  ram[9334]  = 1;
  ram[9335]  = 0;
  ram[9336]  = 0;
  ram[9337]  = 1;
  ram[9338]  = 1;
  ram[9339]  = 1;
  ram[9340]  = 1;
  ram[9341]  = 0;
  ram[9342]  = 1;
  ram[9343]  = 1;
  ram[9344]  = 1;
  ram[9345]  = 1;
  ram[9346]  = 0;
  ram[9347]  = 0;
  ram[9348]  = 1;
  ram[9349]  = 1;
  ram[9350]  = 1;
  ram[9351]  = 1;
  ram[9352]  = 1;
  ram[9353]  = 1;
  ram[9354]  = 1;
  ram[9355]  = 1;
  ram[9356]  = 1;
  ram[9357]  = 1;
  ram[9358]  = 1;
  ram[9359]  = 1;
  ram[9360]  = 1;
  ram[9361]  = 1;
  ram[9362]  = 1;
  ram[9363]  = 1;
  ram[9364]  = 1;
  ram[9365]  = 1;
  ram[9366]  = 1;
  ram[9367]  = 1;
  ram[9368]  = 1;
  ram[9369]  = 0;
  ram[9370]  = 0;
  ram[9371]  = 1;
  ram[9372]  = 1;
  ram[9373]  = 1;
  ram[9374]  = 1;
  ram[9375]  = 1;
  ram[9376]  = 1;
  ram[9377]  = 1;
  ram[9378]  = 1;
  ram[9379]  = 1;
  ram[9380]  = 1;
  ram[9381]  = 1;
  ram[9382]  = 1;
  ram[9383]  = 1;
  ram[9384]  = 1;
  ram[9385]  = 1;
  ram[9386]  = 1;
  ram[9387]  = 1;
  ram[9388]  = 1;
  ram[9389]  = 1;
  ram[9390]  = 1;
  ram[9391]  = 1;
  ram[9392]  = 1;
  ram[9393]  = 1;
  ram[9394]  = 1;
  ram[9395]  = 1;
  ram[9396]  = 1;
  ram[9397]  = 1;
  ram[9398]  = 1;
  ram[9399]  = 1;
  ram[9400]  = 1;
  ram[9401]  = 1;
  ram[9402]  = 1;
  ram[9403]  = 1;
  ram[9404]  = 1;
  ram[9405]  = 1;
  ram[9406]  = 1;
  ram[9407]  = 1;
  ram[9408]  = 1;
  ram[9409]  = 1;
  ram[9410]  = 1;
  ram[9411]  = 1;
  ram[9412]  = 1;
  ram[9413]  = 1;
  ram[9414]  = 1;
  ram[9415]  = 1;
  ram[9416]  = 1;
  ram[9417]  = 1;
  ram[9418]  = 1;
  ram[9419]  = 1;
  ram[9420]  = 0;
  ram[9421]  = 0;
  ram[9422]  = 1;
  ram[9423]  = 1;
  ram[9424]  = 1;
  ram[9425]  = 1;
  ram[9426]  = 0;
  ram[9427]  = 0;
  ram[9428]  = 1;
  ram[9429]  = 1;
  ram[9430]  = 1;
  ram[9431]  = 1;
  ram[9432]  = 1;
  ram[9433]  = 1;
  ram[9434]  = 1;
  ram[9435]  = 0;
  ram[9436]  = 1;
  ram[9437]  = 1;
  ram[9438]  = 1;
  ram[9439]  = 1;
  ram[9440]  = 1;
  ram[9441]  = 1;
  ram[9442]  = 1;
  ram[9443]  = 0;
  ram[9444]  = 0;
  ram[9445]  = 1;
  ram[9446]  = 1;
  ram[9447]  = 1;
  ram[9448]  = 1;
  ram[9449]  = 1;
  ram[9450]  = 0;
  ram[9451]  = 0;
  ram[9452]  = 0;
  ram[9453]  = 1;
  ram[9454]  = 1;
  ram[9455]  = 1;
  ram[9456]  = 1;
  ram[9457]  = 0;
  ram[9458]  = 0;
  ram[9459]  = 1;
  ram[9460]  = 1;
  ram[9461]  = 1;
  ram[9462]  = 1;
  ram[9463]  = 1;
  ram[9464]  = 0;
  ram[9465]  = 0;
  ram[9466]  = 1;
  ram[9467]  = 1;
  ram[9468]  = 1;
  ram[9469]  = 1;
  ram[9470]  = 0;
  ram[9471]  = 0;
  ram[9472]  = 0;
  ram[9473]  = 0;
  ram[9474]  = 0;
  ram[9475]  = 0;
  ram[9476]  = 1;
  ram[9477]  = 1;
  ram[9478]  = 1;
  ram[9479]  = 1;
  ram[9480]  = 1;
  ram[9481]  = 0;
  ram[9482]  = 0;
  ram[9483]  = 1;
  ram[9484]  = 1;
  ram[9485]  = 1;
  ram[9486]  = 1;
  ram[9487]  = 1;
  ram[9488]  = 1;
  ram[9489]  = 1;
  ram[9490]  = 1;
  ram[9491]  = 1;
  ram[9492]  = 1;
  ram[9493]  = 1;
  ram[9494]  = 1;
  ram[9495]  = 1;
  ram[9496]  = 1;
  ram[9497]  = 1;
  ram[9498]  = 1;
  ram[9499]  = 1;
  ram[9500]  = 1;
  ram[9501]  = 1;
  ram[9502]  = 1;
  ram[9503]  = 1;
  ram[9504]  = 1;
  ram[9505]  = 1;
  ram[9506]  = 1;
  ram[9507]  = 1;
  ram[9508]  = 1;
  ram[9509]  = 1;
  ram[9510]  = 1;
  ram[9511]  = 1;
  ram[9512]  = 1;
  ram[9513]  = 1;
  ram[9514]  = 1;
  ram[9515]  = 0;
  ram[9516]  = 0;
  ram[9517]  = 0;
  ram[9518]  = 1;
  ram[9519]  = 1;
  ram[9520]  = 0;
  ram[9521]  = 0;
  ram[9522]  = 0;
  ram[9523]  = 1;
  ram[9524]  = 1;
  ram[9525]  = 1;
  ram[9526]  = 1;
  ram[9527]  = 1;
  ram[9528]  = 0;
  ram[9529]  = 0;
  ram[9530]  = 1;
  ram[9531]  = 1;
  ram[9532]  = 1;
  ram[9533]  = 1;
  ram[9534]  = 1;
  ram[9535]  = 0;
  ram[9536]  = 0;
  ram[9537]  = 1;
  ram[9538]  = 1;
  ram[9539]  = 1;
  ram[9540]  = 1;
  ram[9541]  = 0;
  ram[9542]  = 1;
  ram[9543]  = 1;
  ram[9544]  = 1;
  ram[9545]  = 1;
  ram[9546]  = 0;
  ram[9547]  = 0;
  ram[9548]  = 1;
  ram[9549]  = 1;
  ram[9550]  = 1;
  ram[9551]  = 1;
  ram[9552]  = 1;
  ram[9553]  = 1;
  ram[9554]  = 1;
  ram[9555]  = 1;
  ram[9556]  = 1;
  ram[9557]  = 1;
  ram[9558]  = 1;
  ram[9559]  = 1;
  ram[9560]  = 1;
  ram[9561]  = 1;
  ram[9562]  = 1;
  ram[9563]  = 1;
  ram[9564]  = 1;
  ram[9565]  = 1;
  ram[9566]  = 1;
  ram[9567]  = 1;
  ram[9568]  = 1;
  ram[9569]  = 0;
  ram[9570]  = 0;
  ram[9571]  = 1;
  ram[9572]  = 1;
  ram[9573]  = 1;
  ram[9574]  = 1;
  ram[9575]  = 1;
  ram[9576]  = 1;
  ram[9577]  = 1;
  ram[9578]  = 1;
  ram[9579]  = 1;
  ram[9580]  = 1;
  ram[9581]  = 1;
  ram[9582]  = 1;
  ram[9583]  = 1;
  ram[9584]  = 1;
  ram[9585]  = 1;
  ram[9586]  = 1;
  ram[9587]  = 1;
  ram[9588]  = 1;
  ram[9589]  = 1;
  ram[9590]  = 1;
  ram[9591]  = 1;
  ram[9592]  = 1;
  ram[9593]  = 1;
  ram[9594]  = 1;
  ram[9595]  = 1;
  ram[9596]  = 1;
  ram[9597]  = 1;
  ram[9598]  = 1;
  ram[9599]  = 1;
  ram[9600]  = 1;
  ram[9601]  = 1;
  ram[9602]  = 1;
  ram[9603]  = 1;
  ram[9604]  = 1;
  ram[9605]  = 1;
  ram[9606]  = 1;
  ram[9607]  = 1;
  ram[9608]  = 1;
  ram[9609]  = 1;
  ram[9610]  = 1;
  ram[9611]  = 1;
  ram[9612]  = 1;
  ram[9613]  = 1;
  ram[9614]  = 1;
  ram[9615]  = 1;
  ram[9616]  = 1;
  ram[9617]  = 1;
  ram[9618]  = 1;
  ram[9619]  = 1;
  ram[9620]  = 0;
  ram[9621]  = 0;
  ram[9622]  = 1;
  ram[9623]  = 1;
  ram[9624]  = 1;
  ram[9625]  = 1;
  ram[9626]  = 0;
  ram[9627]  = 0;
  ram[9628]  = 1;
  ram[9629]  = 1;
  ram[9630]  = 1;
  ram[9631]  = 1;
  ram[9632]  = 1;
  ram[9633]  = 1;
  ram[9634]  = 1;
  ram[9635]  = 0;
  ram[9636]  = 1;
  ram[9637]  = 1;
  ram[9638]  = 1;
  ram[9639]  = 1;
  ram[9640]  = 1;
  ram[9641]  = 1;
  ram[9642]  = 1;
  ram[9643]  = 0;
  ram[9644]  = 0;
  ram[9645]  = 1;
  ram[9646]  = 1;
  ram[9647]  = 1;
  ram[9648]  = 1;
  ram[9649]  = 1;
  ram[9650]  = 0;
  ram[9651]  = 0;
  ram[9652]  = 1;
  ram[9653]  = 1;
  ram[9654]  = 1;
  ram[9655]  = 1;
  ram[9656]  = 1;
  ram[9657]  = 0;
  ram[9658]  = 0;
  ram[9659]  = 1;
  ram[9660]  = 1;
  ram[9661]  = 1;
  ram[9662]  = 1;
  ram[9663]  = 1;
  ram[9664]  = 0;
  ram[9665]  = 0;
  ram[9666]  = 1;
  ram[9667]  = 0;
  ram[9668]  = 0;
  ram[9669]  = 0;
  ram[9670]  = 0;
  ram[9671]  = 0;
  ram[9672]  = 0;
  ram[9673]  = 0;
  ram[9674]  = 1;
  ram[9675]  = 1;
  ram[9676]  = 1;
  ram[9677]  = 1;
  ram[9678]  = 1;
  ram[9679]  = 1;
  ram[9680]  = 1;
  ram[9681]  = 0;
  ram[9682]  = 0;
  ram[9683]  = 1;
  ram[9684]  = 1;
  ram[9685]  = 1;
  ram[9686]  = 1;
  ram[9687]  = 1;
  ram[9688]  = 1;
  ram[9689]  = 1;
  ram[9690]  = 1;
  ram[9691]  = 1;
  ram[9692]  = 1;
  ram[9693]  = 1;
  ram[9694]  = 1;
  ram[9695]  = 1;
  ram[9696]  = 1;
  ram[9697]  = 1;
  ram[9698]  = 1;
  ram[9699]  = 1;
  ram[9700]  = 1;
  ram[9701]  = 1;
  ram[9702]  = 1;
  ram[9703]  = 1;
  ram[9704]  = 1;
  ram[9705]  = 1;
  ram[9706]  = 1;
  ram[9707]  = 1;
  ram[9708]  = 1;
  ram[9709]  = 1;
  ram[9710]  = 1;
  ram[9711]  = 1;
  ram[9712]  = 1;
  ram[9713]  = 1;
  ram[9714]  = 1;
  ram[9715]  = 0;
  ram[9716]  = 0;
  ram[9717]  = 0;
  ram[9718]  = 0;
  ram[9719]  = 0;
  ram[9720]  = 0;
  ram[9721]  = 0;
  ram[9722]  = 0;
  ram[9723]  = 0;
  ram[9724]  = 0;
  ram[9725]  = 0;
  ram[9726]  = 1;
  ram[9727]  = 1;
  ram[9728]  = 0;
  ram[9729]  = 0;
  ram[9730]  = 1;
  ram[9731]  = 1;
  ram[9732]  = 1;
  ram[9733]  = 1;
  ram[9734]  = 1;
  ram[9735]  = 0;
  ram[9736]  = 0;
  ram[9737]  = 1;
  ram[9738]  = 1;
  ram[9739]  = 1;
  ram[9740]  = 1;
  ram[9741]  = 0;
  ram[9742]  = 1;
  ram[9743]  = 1;
  ram[9744]  = 1;
  ram[9745]  = 1;
  ram[9746]  = 0;
  ram[9747]  = 0;
  ram[9748]  = 1;
  ram[9749]  = 1;
  ram[9750]  = 1;
  ram[9751]  = 1;
  ram[9752]  = 1;
  ram[9753]  = 1;
  ram[9754]  = 1;
  ram[9755]  = 1;
  ram[9756]  = 1;
  ram[9757]  = 1;
  ram[9758]  = 1;
  ram[9759]  = 1;
  ram[9760]  = 1;
  ram[9761]  = 1;
  ram[9762]  = 1;
  ram[9763]  = 1;
  ram[9764]  = 1;
  ram[9765]  = 1;
  ram[9766]  = 1;
  ram[9767]  = 1;
  ram[9768]  = 1;
  ram[9769]  = 0;
  ram[9770]  = 0;
  ram[9771]  = 1;
  ram[9772]  = 1;
  ram[9773]  = 1;
  ram[9774]  = 1;
  ram[9775]  = 1;
  ram[9776]  = 1;
  ram[9777]  = 1;
  ram[9778]  = 1;
  ram[9779]  = 1;
  ram[9780]  = 1;
  ram[9781]  = 1;
  ram[9782]  = 1;
  ram[9783]  = 1;
  ram[9784]  = 1;
  ram[9785]  = 1;
  ram[9786]  = 1;
  ram[9787]  = 1;
  ram[9788]  = 1;
  ram[9789]  = 1;
  ram[9790]  = 1;
  ram[9791]  = 1;
  ram[9792]  = 1;
  ram[9793]  = 1;
  ram[9794]  = 1;
  ram[9795]  = 1;
  ram[9796]  = 1;
  ram[9797]  = 1;
  ram[9798]  = 1;
  ram[9799]  = 1;
  ram[9800]  = 1;
  ram[9801]  = 1;
  ram[9802]  = 1;
  ram[9803]  = 1;
  ram[9804]  = 1;
  ram[9805]  = 1;
  ram[9806]  = 1;
  ram[9807]  = 1;
  ram[9808]  = 1;
  ram[9809]  = 1;
  ram[9810]  = 1;
  ram[9811]  = 1;
  ram[9812]  = 1;
  ram[9813]  = 1;
  ram[9814]  = 1;
  ram[9815]  = 1;
  ram[9816]  = 1;
  ram[9817]  = 1;
  ram[9818]  = 1;
  ram[9819]  = 1;
  ram[9820]  = 0;
  ram[9821]  = 0;
  ram[9822]  = 1;
  ram[9823]  = 1;
  ram[9824]  = 1;
  ram[9825]  = 1;
  ram[9826]  = 0;
  ram[9827]  = 0;
  ram[9828]  = 1;
  ram[9829]  = 1;
  ram[9830]  = 1;
  ram[9831]  = 1;
  ram[9832]  = 1;
  ram[9833]  = 1;
  ram[9834]  = 1;
  ram[9835]  = 0;
  ram[9836]  = 0;
  ram[9837]  = 0;
  ram[9838]  = 0;
  ram[9839]  = 0;
  ram[9840]  = 0;
  ram[9841]  = 1;
  ram[9842]  = 1;
  ram[9843]  = 1;
  ram[9844]  = 0;
  ram[9845]  = 1;
  ram[9846]  = 1;
  ram[9847]  = 1;
  ram[9848]  = 1;
  ram[9849]  = 0;
  ram[9850]  = 0;
  ram[9851]  = 0;
  ram[9852]  = 1;
  ram[9853]  = 1;
  ram[9854]  = 1;
  ram[9855]  = 1;
  ram[9856]  = 1;
  ram[9857]  = 0;
  ram[9858]  = 0;
  ram[9859]  = 1;
  ram[9860]  = 1;
  ram[9861]  = 1;
  ram[9862]  = 1;
  ram[9863]  = 1;
  ram[9864]  = 0;
  ram[9865]  = 0;
  ram[9866]  = 1;
  ram[9867]  = 0;
  ram[9868]  = 0;
  ram[9869]  = 0;
  ram[9870]  = 0;
  ram[9871]  = 1;
  ram[9872]  = 0;
  ram[9873]  = 0;
  ram[9874]  = 1;
  ram[9875]  = 1;
  ram[9876]  = 1;
  ram[9877]  = 1;
  ram[9878]  = 1;
  ram[9879]  = 1;
  ram[9880]  = 1;
  ram[9881]  = 0;
  ram[9882]  = 0;
  ram[9883]  = 1;
  ram[9884]  = 1;
  ram[9885]  = 1;
  ram[9886]  = 1;
  ram[9887]  = 1;
  ram[9888]  = 1;
  ram[9889]  = 1;
  ram[9890]  = 1;
  ram[9891]  = 1;
  ram[9892]  = 1;
  ram[9893]  = 1;
  ram[9894]  = 1;
  ram[9895]  = 1;
  ram[9896]  = 1;
  ram[9897]  = 1;
  ram[9898]  = 1;
  ram[9899]  = 1;
  ram[9900]  = 1;
  ram[9901]  = 1;
  ram[9902]  = 1;
  ram[9903]  = 1;
  ram[9904]  = 1;
  ram[9905]  = 1;
  ram[9906]  = 1;
  ram[9907]  = 1;
  ram[9908]  = 1;
  ram[9909]  = 1;
  ram[9910]  = 1;
  ram[9911]  = 1;
  ram[9912]  = 1;
  ram[9913]  = 1;
  ram[9914]  = 1;
  ram[9915]  = 1;
  ram[9916]  = 1;
  ram[9917]  = 1;
  ram[9918]  = 1;
  ram[9919]  = 1;
  ram[9920]  = 1;
  ram[9921]  = 0;
  ram[9922]  = 0;
  ram[9923]  = 1;
  ram[9924]  = 1;
  ram[9925]  = 1;
  ram[9926]  = 1;
  ram[9927]  = 1;
  ram[9928]  = 0;
  ram[9929]  = 0;
  ram[9930]  = 1;
  ram[9931]  = 1;
  ram[9932]  = 1;
  ram[9933]  = 1;
  ram[9934]  = 1;
  ram[9935]  = 0;
  ram[9936]  = 0;
  ram[9937]  = 1;
  ram[9938]  = 1;
  ram[9939]  = 1;
  ram[9940]  = 1;
  ram[9941]  = 0;
  ram[9942]  = 1;
  ram[9943]  = 1;
  ram[9944]  = 1;
  ram[9945]  = 1;
  ram[9946]  = 0;
  ram[9947]  = 0;
  ram[9948]  = 1;
  ram[9949]  = 1;
  ram[9950]  = 1;
  ram[9951]  = 1;
  ram[9952]  = 1;
  ram[9953]  = 1;
  ram[9954]  = 1;
  ram[9955]  = 1;
  ram[9956]  = 1;
  ram[9957]  = 1;
  ram[9958]  = 1;
  ram[9959]  = 1;
  ram[9960]  = 1;
  ram[9961]  = 1;
  ram[9962]  = 1;
  ram[9963]  = 1;
  ram[9964]  = 1;
  ram[9965]  = 1;
  ram[9966]  = 1;
  ram[9967]  = 1;
  ram[9968]  = 1;
  ram[9969]  = 0;
  ram[9970]  = 0;
  ram[9971]  = 1;
  ram[9972]  = 1;
  ram[9973]  = 1;
  ram[9974]  = 1;
  ram[9975]  = 1;
  ram[9976]  = 1;
  ram[9977]  = 1;
  ram[9978]  = 1;
  ram[9979]  = 1;
  ram[9980]  = 1;
  ram[9981]  = 1;
  ram[9982]  = 1;
  ram[9983]  = 1;
  ram[9984]  = 1;
  ram[9985]  = 1;
  ram[9986]  = 1;
  ram[9987]  = 1;
  ram[9988]  = 1;
  ram[9989]  = 1;
  ram[9990]  = 1;
  ram[9991]  = 1;
  ram[9992]  = 1;
  ram[9993]  = 1;
  ram[9994]  = 1;
  ram[9995]  = 1;
  ram[9996]  = 1;
  ram[9997]  = 1;
  ram[9998]  = 1;
  ram[9999]  = 1;
  ram[10000]  = 1;
  ram[10001]  = 1;
  ram[10002]  = 1;
  ram[10003]  = 1;
  ram[10004]  = 1;
  ram[10005]  = 1;
  ram[10006]  = 1;
  ram[10007]  = 1;
  ram[10008]  = 1;
  ram[10009]  = 1;
  ram[10010]  = 1;
  ram[10011]  = 1;
  ram[10012]  = 1;
  ram[10013]  = 1;
  ram[10014]  = 1;
  ram[10015]  = 1;
  ram[10016]  = 1;
  ram[10017]  = 1;
  ram[10018]  = 1;
  ram[10019]  = 1;
  ram[10020]  = 0;
  ram[10021]  = 0;
  ram[10022]  = 1;
  ram[10023]  = 1;
  ram[10024]  = 1;
  ram[10025]  = 1;
  ram[10026]  = 0;
  ram[10027]  = 0;
  ram[10028]  = 1;
  ram[10029]  = 1;
  ram[10030]  = 1;
  ram[10031]  = 1;
  ram[10032]  = 1;
  ram[10033]  = 0;
  ram[10034]  = 0;
  ram[10035]  = 0;
  ram[10036]  = 0;
  ram[10037]  = 0;
  ram[10038]  = 0;
  ram[10039]  = 0;
  ram[10040]  = 0;
  ram[10041]  = 1;
  ram[10042]  = 1;
  ram[10043]  = 1;
  ram[10044]  = 0;
  ram[10045]  = 1;
  ram[10046]  = 1;
  ram[10047]  = 1;
  ram[10048]  = 0;
  ram[10049]  = 0;
  ram[10050]  = 0;
  ram[10051]  = 1;
  ram[10052]  = 1;
  ram[10053]  = 1;
  ram[10054]  = 1;
  ram[10055]  = 1;
  ram[10056]  = 1;
  ram[10057]  = 0;
  ram[10058]  = 0;
  ram[10059]  = 1;
  ram[10060]  = 1;
  ram[10061]  = 1;
  ram[10062]  = 1;
  ram[10063]  = 1;
  ram[10064]  = 0;
  ram[10065]  = 0;
  ram[10066]  = 1;
  ram[10067]  = 1;
  ram[10068]  = 0;
  ram[10069]  = 1;
  ram[10070]  = 1;
  ram[10071]  = 1;
  ram[10072]  = 0;
  ram[10073]  = 0;
  ram[10074]  = 1;
  ram[10075]  = 1;
  ram[10076]  = 1;
  ram[10077]  = 1;
  ram[10078]  = 1;
  ram[10079]  = 1;
  ram[10080]  = 1;
  ram[10081]  = 0;
  ram[10082]  = 0;
  ram[10083]  = 1;
  ram[10084]  = 1;
  ram[10085]  = 1;
  ram[10086]  = 1;
  ram[10087]  = 1;
  ram[10088]  = 1;
  ram[10089]  = 1;
  ram[10090]  = 1;
  ram[10091]  = 1;
  ram[10092]  = 1;
  ram[10093]  = 1;
  ram[10094]  = 1;
  ram[10095]  = 1;
  ram[10096]  = 1;
  ram[10097]  = 1;
  ram[10098]  = 1;
  ram[10099]  = 1;
  ram[10100]  = 1;
  ram[10101]  = 1;
  ram[10102]  = 1;
  ram[10103]  = 1;
  ram[10104]  = 1;
  ram[10105]  = 1;
  ram[10106]  = 1;
  ram[10107]  = 1;
  ram[10108]  = 1;
  ram[10109]  = 1;
  ram[10110]  = 1;
  ram[10111]  = 1;
  ram[10112]  = 1;
  ram[10113]  = 1;
  ram[10114]  = 1;
  ram[10115]  = 1;
  ram[10116]  = 1;
  ram[10117]  = 1;
  ram[10118]  = 1;
  ram[10119]  = 1;
  ram[10120]  = 1;
  ram[10121]  = 0;
  ram[10122]  = 0;
  ram[10123]  = 1;
  ram[10124]  = 1;
  ram[10125]  = 1;
  ram[10126]  = 1;
  ram[10127]  = 1;
  ram[10128]  = 0;
  ram[10129]  = 0;
  ram[10130]  = 0;
  ram[10131]  = 0;
  ram[10132]  = 0;
  ram[10133]  = 0;
  ram[10134]  = 0;
  ram[10135]  = 0;
  ram[10136]  = 0;
  ram[10137]  = 1;
  ram[10138]  = 1;
  ram[10139]  = 1;
  ram[10140]  = 1;
  ram[10141]  = 0;
  ram[10142]  = 1;
  ram[10143]  = 1;
  ram[10144]  = 1;
  ram[10145]  = 1;
  ram[10146]  = 0;
  ram[10147]  = 0;
  ram[10148]  = 1;
  ram[10149]  = 1;
  ram[10150]  = 1;
  ram[10151]  = 1;
  ram[10152]  = 1;
  ram[10153]  = 1;
  ram[10154]  = 1;
  ram[10155]  = 1;
  ram[10156]  = 1;
  ram[10157]  = 1;
  ram[10158]  = 1;
  ram[10159]  = 1;
  ram[10160]  = 1;
  ram[10161]  = 1;
  ram[10162]  = 1;
  ram[10163]  = 1;
  ram[10164]  = 1;
  ram[10165]  = 1;
  ram[10166]  = 1;
  ram[10167]  = 1;
  ram[10168]  = 1;
  ram[10169]  = 0;
  ram[10170]  = 0;
  ram[10171]  = 1;
  ram[10172]  = 1;
  ram[10173]  = 1;
  ram[10174]  = 1;
  ram[10175]  = 1;
  ram[10176]  = 1;
  ram[10177]  = 1;
  ram[10178]  = 1;
  ram[10179]  = 1;
  ram[10180]  = 1;
  ram[10181]  = 1;
  ram[10182]  = 1;
  ram[10183]  = 1;
  ram[10184]  = 1;
  ram[10185]  = 1;
  ram[10186]  = 1;
  ram[10187]  = 1;
  ram[10188]  = 1;
  ram[10189]  = 1;
  ram[10190]  = 1;
  ram[10191]  = 1;
  ram[10192]  = 1;
  ram[10193]  = 1;
  ram[10194]  = 1;
  ram[10195]  = 1;
  ram[10196]  = 1;
  ram[10197]  = 1;
  ram[10198]  = 1;
  ram[10199]  = 1;
  ram[10200]  = 1;
  ram[10201]  = 1;
  ram[10202]  = 1;
  ram[10203]  = 1;
  ram[10204]  = 1;
  ram[10205]  = 1;
  ram[10206]  = 1;
  ram[10207]  = 1;
  ram[10208]  = 1;
  ram[10209]  = 1;
  ram[10210]  = 1;
  ram[10211]  = 1;
  ram[10212]  = 1;
  ram[10213]  = 1;
  ram[10214]  = 1;
  ram[10215]  = 1;
  ram[10216]  = 1;
  ram[10217]  = 1;
  ram[10218]  = 1;
  ram[10219]  = 1;
  ram[10220]  = 0;
  ram[10221]  = 0;
  ram[10222]  = 1;
  ram[10223]  = 1;
  ram[10224]  = 1;
  ram[10225]  = 1;
  ram[10226]  = 0;
  ram[10227]  = 0;
  ram[10228]  = 1;
  ram[10229]  = 0;
  ram[10230]  = 0;
  ram[10231]  = 0;
  ram[10232]  = 0;
  ram[10233]  = 0;
  ram[10234]  = 0;
  ram[10235]  = 0;
  ram[10236]  = 0;
  ram[10237]  = 1;
  ram[10238]  = 1;
  ram[10239]  = 1;
  ram[10240]  = 1;
  ram[10241]  = 1;
  ram[10242]  = 1;
  ram[10243]  = 1;
  ram[10244]  = 0;
  ram[10245]  = 0;
  ram[10246]  = 1;
  ram[10247]  = 1;
  ram[10248]  = 0;
  ram[10249]  = 0;
  ram[10250]  = 1;
  ram[10251]  = 1;
  ram[10252]  = 1;
  ram[10253]  = 1;
  ram[10254]  = 1;
  ram[10255]  = 1;
  ram[10256]  = 1;
  ram[10257]  = 0;
  ram[10258]  = 0;
  ram[10259]  = 1;
  ram[10260]  = 1;
  ram[10261]  = 1;
  ram[10262]  = 1;
  ram[10263]  = 1;
  ram[10264]  = 0;
  ram[10265]  = 0;
  ram[10266]  = 1;
  ram[10267]  = 1;
  ram[10268]  = 1;
  ram[10269]  = 1;
  ram[10270]  = 1;
  ram[10271]  = 1;
  ram[10272]  = 0;
  ram[10273]  = 0;
  ram[10274]  = 1;
  ram[10275]  = 1;
  ram[10276]  = 1;
  ram[10277]  = 1;
  ram[10278]  = 1;
  ram[10279]  = 1;
  ram[10280]  = 1;
  ram[10281]  = 0;
  ram[10282]  = 0;
  ram[10283]  = 1;
  ram[10284]  = 1;
  ram[10285]  = 1;
  ram[10286]  = 1;
  ram[10287]  = 1;
  ram[10288]  = 1;
  ram[10289]  = 1;
  ram[10290]  = 1;
  ram[10291]  = 1;
  ram[10292]  = 1;
  ram[10293]  = 1;
  ram[10294]  = 1;
  ram[10295]  = 1;
  ram[10296]  = 1;
  ram[10297]  = 1;
  ram[10298]  = 1;
  ram[10299]  = 1;
  ram[10300]  = 1;
  ram[10301]  = 1;
  ram[10302]  = 1;
  ram[10303]  = 1;
  ram[10304]  = 1;
  ram[10305]  = 1;
  ram[10306]  = 1;
  ram[10307]  = 1;
  ram[10308]  = 1;
  ram[10309]  = 1;
  ram[10310]  = 1;
  ram[10311]  = 1;
  ram[10312]  = 1;
  ram[10313]  = 1;
  ram[10314]  = 1;
  ram[10315]  = 1;
  ram[10316]  = 1;
  ram[10317]  = 1;
  ram[10318]  = 1;
  ram[10319]  = 1;
  ram[10320]  = 1;
  ram[10321]  = 0;
  ram[10322]  = 0;
  ram[10323]  = 1;
  ram[10324]  = 1;
  ram[10325]  = 1;
  ram[10326]  = 1;
  ram[10327]  = 1;
  ram[10328]  = 0;
  ram[10329]  = 0;
  ram[10330]  = 1;
  ram[10331]  = 1;
  ram[10332]  = 1;
  ram[10333]  = 1;
  ram[10334]  = 1;
  ram[10335]  = 0;
  ram[10336]  = 0;
  ram[10337]  = 1;
  ram[10338]  = 1;
  ram[10339]  = 1;
  ram[10340]  = 1;
  ram[10341]  = 0;
  ram[10342]  = 1;
  ram[10343]  = 1;
  ram[10344]  = 1;
  ram[10345]  = 1;
  ram[10346]  = 0;
  ram[10347]  = 0;
  ram[10348]  = 1;
  ram[10349]  = 1;
  ram[10350]  = 1;
  ram[10351]  = 1;
  ram[10352]  = 1;
  ram[10353]  = 1;
  ram[10354]  = 1;
  ram[10355]  = 1;
  ram[10356]  = 1;
  ram[10357]  = 1;
  ram[10358]  = 1;
  ram[10359]  = 1;
  ram[10360]  = 1;
  ram[10361]  = 1;
  ram[10362]  = 1;
  ram[10363]  = 1;
  ram[10364]  = 1;
  ram[10365]  = 1;
  ram[10366]  = 1;
  ram[10367]  = 1;
  ram[10368]  = 1;
  ram[10369]  = 0;
  ram[10370]  = 0;
  ram[10371]  = 1;
  ram[10372]  = 1;
  ram[10373]  = 1;
  ram[10374]  = 1;
  ram[10375]  = 1;
  ram[10376]  = 1;
  ram[10377]  = 1;
  ram[10378]  = 1;
  ram[10379]  = 1;
  ram[10380]  = 1;
  ram[10381]  = 1;
  ram[10382]  = 1;
  ram[10383]  = 1;
  ram[10384]  = 1;
  ram[10385]  = 1;
  ram[10386]  = 1;
  ram[10387]  = 1;
  ram[10388]  = 1;
  ram[10389]  = 1;
  ram[10390]  = 1;
  ram[10391]  = 1;
  ram[10392]  = 1;
  ram[10393]  = 1;
  ram[10394]  = 1;
  ram[10395]  = 1;
  ram[10396]  = 1;
  ram[10397]  = 1;
  ram[10398]  = 1;
  ram[10399]  = 1;
  ram[10400]  = 1;
  ram[10401]  = 1;
  ram[10402]  = 1;
  ram[10403]  = 1;
  ram[10404]  = 1;
  ram[10405]  = 1;
  ram[10406]  = 1;
  ram[10407]  = 1;
  ram[10408]  = 1;
  ram[10409]  = 1;
  ram[10410]  = 1;
  ram[10411]  = 1;
  ram[10412]  = 1;
  ram[10413]  = 1;
  ram[10414]  = 1;
  ram[10415]  = 1;
  ram[10416]  = 1;
  ram[10417]  = 1;
  ram[10418]  = 1;
  ram[10419]  = 1;
  ram[10420]  = 0;
  ram[10421]  = 0;
  ram[10422]  = 1;
  ram[10423]  = 1;
  ram[10424]  = 1;
  ram[10425]  = 1;
  ram[10426]  = 0;
  ram[10427]  = 0;
  ram[10428]  = 1;
  ram[10429]  = 1;
  ram[10430]  = 0;
  ram[10431]  = 0;
  ram[10432]  = 0;
  ram[10433]  = 0;
  ram[10434]  = 0;
  ram[10435]  = 0;
  ram[10436]  = 1;
  ram[10437]  = 1;
  ram[10438]  = 1;
  ram[10439]  = 1;
  ram[10440]  = 1;
  ram[10441]  = 1;
  ram[10442]  = 1;
  ram[10443]  = 1;
  ram[10444]  = 0;
  ram[10445]  = 0;
  ram[10446]  = 1;
  ram[10447]  = 0;
  ram[10448]  = 0;
  ram[10449]  = 1;
  ram[10450]  = 1;
  ram[10451]  = 1;
  ram[10452]  = 1;
  ram[10453]  = 1;
  ram[10454]  = 1;
  ram[10455]  = 1;
  ram[10456]  = 1;
  ram[10457]  = 0;
  ram[10458]  = 0;
  ram[10459]  = 1;
  ram[10460]  = 1;
  ram[10461]  = 1;
  ram[10462]  = 1;
  ram[10463]  = 1;
  ram[10464]  = 0;
  ram[10465]  = 0;
  ram[10466]  = 1;
  ram[10467]  = 1;
  ram[10468]  = 1;
  ram[10469]  = 1;
  ram[10470]  = 1;
  ram[10471]  = 1;
  ram[10472]  = 0;
  ram[10473]  = 0;
  ram[10474]  = 1;
  ram[10475]  = 1;
  ram[10476]  = 1;
  ram[10477]  = 1;
  ram[10478]  = 1;
  ram[10479]  = 1;
  ram[10480]  = 1;
  ram[10481]  = 0;
  ram[10482]  = 0;
  ram[10483]  = 1;
  ram[10484]  = 1;
  ram[10485]  = 1;
  ram[10486]  = 1;
  ram[10487]  = 1;
  ram[10488]  = 1;
  ram[10489]  = 1;
  ram[10490]  = 1;
  ram[10491]  = 1;
  ram[10492]  = 1;
  ram[10493]  = 1;
  ram[10494]  = 1;
  ram[10495]  = 1;
  ram[10496]  = 1;
  ram[10497]  = 1;
  ram[10498]  = 1;
  ram[10499]  = 1;
  ram[10500]  = 1;
  ram[10501]  = 1;
  ram[10502]  = 1;
  ram[10503]  = 1;
  ram[10504]  = 1;
  ram[10505]  = 1;
  ram[10506]  = 1;
  ram[10507]  = 1;
  ram[10508]  = 1;
  ram[10509]  = 1;
  ram[10510]  = 1;
  ram[10511]  = 1;
  ram[10512]  = 1;
  ram[10513]  = 1;
  ram[10514]  = 1;
  ram[10515]  = 1;
  ram[10516]  = 1;
  ram[10517]  = 1;
  ram[10518]  = 1;
  ram[10519]  = 1;
  ram[10520]  = 1;
  ram[10521]  = 0;
  ram[10522]  = 0;
  ram[10523]  = 1;
  ram[10524]  = 1;
  ram[10525]  = 1;
  ram[10526]  = 1;
  ram[10527]  = 1;
  ram[10528]  = 0;
  ram[10529]  = 0;
  ram[10530]  = 1;
  ram[10531]  = 1;
  ram[10532]  = 1;
  ram[10533]  = 1;
  ram[10534]  = 1;
  ram[10535]  = 0;
  ram[10536]  = 0;
  ram[10537]  = 1;
  ram[10538]  = 1;
  ram[10539]  = 1;
  ram[10540]  = 1;
  ram[10541]  = 0;
  ram[10542]  = 1;
  ram[10543]  = 1;
  ram[10544]  = 1;
  ram[10545]  = 1;
  ram[10546]  = 0;
  ram[10547]  = 0;
  ram[10548]  = 1;
  ram[10549]  = 1;
  ram[10550]  = 1;
  ram[10551]  = 1;
  ram[10552]  = 1;
  ram[10553]  = 1;
  ram[10554]  = 1;
  ram[10555]  = 1;
  ram[10556]  = 1;
  ram[10557]  = 1;
  ram[10558]  = 1;
  ram[10559]  = 1;
  ram[10560]  = 1;
  ram[10561]  = 1;
  ram[10562]  = 1;
  ram[10563]  = 1;
  ram[10564]  = 1;
  ram[10565]  = 1;
  ram[10566]  = 1;
  ram[10567]  = 1;
  ram[10568]  = 1;
  ram[10569]  = 0;
  ram[10570]  = 0;
  ram[10571]  = 1;
  ram[10572]  = 1;
  ram[10573]  = 1;
  ram[10574]  = 1;
  ram[10575]  = 1;
  ram[10576]  = 1;
  ram[10577]  = 1;
  ram[10578]  = 1;
  ram[10579]  = 1;
  ram[10580]  = 1;
  ram[10581]  = 1;
  ram[10582]  = 1;
  ram[10583]  = 1;
  ram[10584]  = 1;
  ram[10585]  = 1;
  ram[10586]  = 1;
  ram[10587]  = 1;
  ram[10588]  = 1;
  ram[10589]  = 1;
  ram[10590]  = 1;
  ram[10591]  = 1;
  ram[10592]  = 1;
  ram[10593]  = 1;
  ram[10594]  = 1;
  ram[10595]  = 1;
  ram[10596]  = 1;
  ram[10597]  = 1;
  ram[10598]  = 1;
  ram[10599]  = 1;
  ram[10600]  = 1;
  ram[10601]  = 1;
  ram[10602]  = 1;
  ram[10603]  = 1;
  ram[10604]  = 1;
  ram[10605]  = 1;
  ram[10606]  = 1;
  ram[10607]  = 1;
  ram[10608]  = 1;
  ram[10609]  = 1;
  ram[10610]  = 1;
  ram[10611]  = 1;
  ram[10612]  = 1;
  ram[10613]  = 1;
  ram[10614]  = 1;
  ram[10615]  = 1;
  ram[10616]  = 1;
  ram[10617]  = 1;
  ram[10618]  = 1;
  ram[10619]  = 1;
  ram[10620]  = 0;
  ram[10621]  = 0;
  ram[10622]  = 1;
  ram[10623]  = 1;
  ram[10624]  = 1;
  ram[10625]  = 1;
  ram[10626]  = 0;
  ram[10627]  = 0;
  ram[10628]  = 1;
  ram[10629]  = 1;
  ram[10630]  = 1;
  ram[10631]  = 1;
  ram[10632]  = 1;
  ram[10633]  = 1;
  ram[10634]  = 1;
  ram[10635]  = 0;
  ram[10636]  = 1;
  ram[10637]  = 1;
  ram[10638]  = 1;
  ram[10639]  = 1;
  ram[10640]  = 1;
  ram[10641]  = 1;
  ram[10642]  = 1;
  ram[10643]  = 1;
  ram[10644]  = 0;
  ram[10645]  = 0;
  ram[10646]  = 0;
  ram[10647]  = 0;
  ram[10648]  = 0;
  ram[10649]  = 1;
  ram[10650]  = 1;
  ram[10651]  = 1;
  ram[10652]  = 1;
  ram[10653]  = 1;
  ram[10654]  = 1;
  ram[10655]  = 1;
  ram[10656]  = 1;
  ram[10657]  = 0;
  ram[10658]  = 0;
  ram[10659]  = 1;
  ram[10660]  = 1;
  ram[10661]  = 1;
  ram[10662]  = 1;
  ram[10663]  = 1;
  ram[10664]  = 0;
  ram[10665]  = 0;
  ram[10666]  = 1;
  ram[10667]  = 1;
  ram[10668]  = 1;
  ram[10669]  = 1;
  ram[10670]  = 1;
  ram[10671]  = 1;
  ram[10672]  = 0;
  ram[10673]  = 0;
  ram[10674]  = 1;
  ram[10675]  = 1;
  ram[10676]  = 1;
  ram[10677]  = 1;
  ram[10678]  = 1;
  ram[10679]  = 1;
  ram[10680]  = 1;
  ram[10681]  = 0;
  ram[10682]  = 0;
  ram[10683]  = 1;
  ram[10684]  = 1;
  ram[10685]  = 1;
  ram[10686]  = 1;
  ram[10687]  = 1;
  ram[10688]  = 1;
  ram[10689]  = 0;
  ram[10690]  = 0;
  ram[10691]  = 1;
  ram[10692]  = 1;
  ram[10693]  = 1;
  ram[10694]  = 1;
  ram[10695]  = 1;
  ram[10696]  = 1;
  ram[10697]  = 1;
  ram[10698]  = 1;
  ram[10699]  = 1;
  ram[10700]  = 1;
  ram[10701]  = 1;
  ram[10702]  = 1;
  ram[10703]  = 1;
  ram[10704]  = 1;
  ram[10705]  = 1;
  ram[10706]  = 1;
  ram[10707]  = 1;
  ram[10708]  = 1;
  ram[10709]  = 1;
  ram[10710]  = 1;
  ram[10711]  = 1;
  ram[10712]  = 1;
  ram[10713]  = 1;
  ram[10714]  = 1;
  ram[10715]  = 1;
  ram[10716]  = 1;
  ram[10717]  = 1;
  ram[10718]  = 1;
  ram[10719]  = 1;
  ram[10720]  = 1;
  ram[10721]  = 0;
  ram[10722]  = 0;
  ram[10723]  = 1;
  ram[10724]  = 1;
  ram[10725]  = 1;
  ram[10726]  = 1;
  ram[10727]  = 1;
  ram[10728]  = 0;
  ram[10729]  = 0;
  ram[10730]  = 1;
  ram[10731]  = 1;
  ram[10732]  = 1;
  ram[10733]  = 1;
  ram[10734]  = 1;
  ram[10735]  = 0;
  ram[10736]  = 0;
  ram[10737]  = 1;
  ram[10738]  = 1;
  ram[10739]  = 1;
  ram[10740]  = 1;
  ram[10741]  = 0;
  ram[10742]  = 1;
  ram[10743]  = 1;
  ram[10744]  = 1;
  ram[10745]  = 1;
  ram[10746]  = 0;
  ram[10747]  = 0;
  ram[10748]  = 1;
  ram[10749]  = 1;
  ram[10750]  = 1;
  ram[10751]  = 1;
  ram[10752]  = 1;
  ram[10753]  = 1;
  ram[10754]  = 1;
  ram[10755]  = 1;
  ram[10756]  = 1;
  ram[10757]  = 1;
  ram[10758]  = 1;
  ram[10759]  = 1;
  ram[10760]  = 1;
  ram[10761]  = 1;
  ram[10762]  = 1;
  ram[10763]  = 1;
  ram[10764]  = 1;
  ram[10765]  = 1;
  ram[10766]  = 1;
  ram[10767]  = 1;
  ram[10768]  = 1;
  ram[10769]  = 0;
  ram[10770]  = 0;
  ram[10771]  = 1;
  ram[10772]  = 1;
  ram[10773]  = 1;
  ram[10774]  = 1;
  ram[10775]  = 1;
  ram[10776]  = 1;
  ram[10777]  = 1;
  ram[10778]  = 1;
  ram[10779]  = 1;
  ram[10780]  = 1;
  ram[10781]  = 1;
  ram[10782]  = 1;
  ram[10783]  = 1;
  ram[10784]  = 1;
  ram[10785]  = 1;
  ram[10786]  = 1;
  ram[10787]  = 1;
  ram[10788]  = 1;
  ram[10789]  = 1;
  ram[10790]  = 1;
  ram[10791]  = 1;
  ram[10792]  = 1;
  ram[10793]  = 1;
  ram[10794]  = 1;
  ram[10795]  = 1;
  ram[10796]  = 1;
  ram[10797]  = 1;
  ram[10798]  = 1;
  ram[10799]  = 1;
  ram[10800]  = 1;
  ram[10801]  = 1;
  ram[10802]  = 1;
  ram[10803]  = 1;
  ram[10804]  = 1;
  ram[10805]  = 1;
  ram[10806]  = 1;
  ram[10807]  = 1;
  ram[10808]  = 1;
  ram[10809]  = 1;
  ram[10810]  = 1;
  ram[10811]  = 1;
  ram[10812]  = 1;
  ram[10813]  = 1;
  ram[10814]  = 1;
  ram[10815]  = 1;
  ram[10816]  = 1;
  ram[10817]  = 1;
  ram[10818]  = 1;
  ram[10819]  = 1;
  ram[10820]  = 0;
  ram[10821]  = 0;
  ram[10822]  = 1;
  ram[10823]  = 1;
  ram[10824]  = 1;
  ram[10825]  = 1;
  ram[10826]  = 0;
  ram[10827]  = 0;
  ram[10828]  = 1;
  ram[10829]  = 1;
  ram[10830]  = 1;
  ram[10831]  = 1;
  ram[10832]  = 1;
  ram[10833]  = 1;
  ram[10834]  = 1;
  ram[10835]  = 0;
  ram[10836]  = 1;
  ram[10837]  = 1;
  ram[10838]  = 1;
  ram[10839]  = 1;
  ram[10840]  = 1;
  ram[10841]  = 1;
  ram[10842]  = 1;
  ram[10843]  = 1;
  ram[10844]  = 0;
  ram[10845]  = 0;
  ram[10846]  = 0;
  ram[10847]  = 0;
  ram[10848]  = 1;
  ram[10849]  = 1;
  ram[10850]  = 1;
  ram[10851]  = 1;
  ram[10852]  = 1;
  ram[10853]  = 1;
  ram[10854]  = 1;
  ram[10855]  = 1;
  ram[10856]  = 1;
  ram[10857]  = 0;
  ram[10858]  = 0;
  ram[10859]  = 1;
  ram[10860]  = 1;
  ram[10861]  = 1;
  ram[10862]  = 1;
  ram[10863]  = 1;
  ram[10864]  = 0;
  ram[10865]  = 0;
  ram[10866]  = 1;
  ram[10867]  = 1;
  ram[10868]  = 1;
  ram[10869]  = 1;
  ram[10870]  = 1;
  ram[10871]  = 1;
  ram[10872]  = 0;
  ram[10873]  = 0;
  ram[10874]  = 1;
  ram[10875]  = 1;
  ram[10876]  = 1;
  ram[10877]  = 1;
  ram[10878]  = 1;
  ram[10879]  = 1;
  ram[10880]  = 1;
  ram[10881]  = 0;
  ram[10882]  = 0;
  ram[10883]  = 1;
  ram[10884]  = 1;
  ram[10885]  = 1;
  ram[10886]  = 1;
  ram[10887]  = 1;
  ram[10888]  = 1;
  ram[10889]  = 0;
  ram[10890]  = 0;
  ram[10891]  = 1;
  ram[10892]  = 1;
  ram[10893]  = 1;
  ram[10894]  = 1;
  ram[10895]  = 1;
  ram[10896]  = 1;
  ram[10897]  = 1;
  ram[10898]  = 1;
  ram[10899]  = 1;
  ram[10900]  = 1;
  ram[10901]  = 1;
  ram[10902]  = 1;
  ram[10903]  = 1;
  ram[10904]  = 1;
  ram[10905]  = 1;
  ram[10906]  = 1;
  ram[10907]  = 1;
  ram[10908]  = 1;
  ram[10909]  = 1;
  ram[10910]  = 1;
  ram[10911]  = 1;
  ram[10912]  = 1;
  ram[10913]  = 1;
  ram[10914]  = 1;
  ram[10915]  = 1;
  ram[10916]  = 1;
  ram[10917]  = 1;
  ram[10918]  = 1;
  ram[10919]  = 1;
  ram[10920]  = 1;
  ram[10921]  = 0;
  ram[10922]  = 0;
  ram[10923]  = 1;
  ram[10924]  = 1;
  ram[10925]  = 1;
  ram[10926]  = 1;
  ram[10927]  = 1;
  ram[10928]  = 0;
  ram[10929]  = 0;
  ram[10930]  = 1;
  ram[10931]  = 1;
  ram[10932]  = 1;
  ram[10933]  = 1;
  ram[10934]  = 1;
  ram[10935]  = 0;
  ram[10936]  = 0;
  ram[10937]  = 1;
  ram[10938]  = 1;
  ram[10939]  = 1;
  ram[10940]  = 1;
  ram[10941]  = 0;
  ram[10942]  = 1;
  ram[10943]  = 1;
  ram[10944]  = 1;
  ram[10945]  = 1;
  ram[10946]  = 0;
  ram[10947]  = 0;
  ram[10948]  = 1;
  ram[10949]  = 1;
  ram[10950]  = 1;
  ram[10951]  = 1;
  ram[10952]  = 1;
  ram[10953]  = 1;
  ram[10954]  = 1;
  ram[10955]  = 1;
  ram[10956]  = 1;
  ram[10957]  = 1;
  ram[10958]  = 1;
  ram[10959]  = 1;
  ram[10960]  = 1;
  ram[10961]  = 1;
  ram[10962]  = 1;
  ram[10963]  = 1;
  ram[10964]  = 1;
  ram[10965]  = 1;
  ram[10966]  = 1;
  ram[10967]  = 1;
  ram[10968]  = 1;
  ram[10969]  = 0;
  ram[10970]  = 0;
  ram[10971]  = 1;
  ram[10972]  = 1;
  ram[10973]  = 1;
  ram[10974]  = 1;
  ram[10975]  = 1;
  ram[10976]  = 1;
  ram[10977]  = 1;
  ram[10978]  = 1;
  ram[10979]  = 1;
  ram[10980]  = 1;
  ram[10981]  = 1;
  ram[10982]  = 1;
  ram[10983]  = 1;
  ram[10984]  = 1;
  ram[10985]  = 1;
  ram[10986]  = 1;
  ram[10987]  = 1;
  ram[10988]  = 1;
  ram[10989]  = 1;
  ram[10990]  = 1;
  ram[10991]  = 1;
  ram[10992]  = 1;
  ram[10993]  = 1;
  ram[10994]  = 1;
  ram[10995]  = 1;
  ram[10996]  = 1;
  ram[10997]  = 1;
  ram[10998]  = 1;
  ram[10999]  = 1;
  ram[11000]  = 1;
  ram[11001]  = 1;
  ram[11002]  = 1;
  ram[11003]  = 1;
  ram[11004]  = 1;
  ram[11005]  = 1;
  ram[11006]  = 1;
  ram[11007]  = 1;
  ram[11008]  = 1;
  ram[11009]  = 1;
  ram[11010]  = 1;
  ram[11011]  = 1;
  ram[11012]  = 1;
  ram[11013]  = 1;
  ram[11014]  = 1;
  ram[11015]  = 1;
  ram[11016]  = 1;
  ram[11017]  = 1;
  ram[11018]  = 1;
  ram[11019]  = 1;
  ram[11020]  = 0;
  ram[11021]  = 0;
  ram[11022]  = 1;
  ram[11023]  = 1;
  ram[11024]  = 1;
  ram[11025]  = 0;
  ram[11026]  = 0;
  ram[11027]  = 0;
  ram[11028]  = 1;
  ram[11029]  = 1;
  ram[11030]  = 1;
  ram[11031]  = 1;
  ram[11032]  = 1;
  ram[11033]  = 1;
  ram[11034]  = 1;
  ram[11035]  = 0;
  ram[11036]  = 1;
  ram[11037]  = 1;
  ram[11038]  = 1;
  ram[11039]  = 1;
  ram[11040]  = 1;
  ram[11041]  = 1;
  ram[11042]  = 1;
  ram[11043]  = 1;
  ram[11044]  = 0;
  ram[11045]  = 0;
  ram[11046]  = 0;
  ram[11047]  = 1;
  ram[11048]  = 1;
  ram[11049]  = 1;
  ram[11050]  = 1;
  ram[11051]  = 1;
  ram[11052]  = 1;
  ram[11053]  = 1;
  ram[11054]  = 1;
  ram[11055]  = 1;
  ram[11056]  = 1;
  ram[11057]  = 0;
  ram[11058]  = 0;
  ram[11059]  = 0;
  ram[11060]  = 0;
  ram[11061]  = 0;
  ram[11062]  = 0;
  ram[11063]  = 0;
  ram[11064]  = 0;
  ram[11065]  = 0;
  ram[11066]  = 1;
  ram[11067]  = 1;
  ram[11068]  = 1;
  ram[11069]  = 1;
  ram[11070]  = 1;
  ram[11071]  = 1;
  ram[11072]  = 0;
  ram[11073]  = 0;
  ram[11074]  = 1;
  ram[11075]  = 1;
  ram[11076]  = 1;
  ram[11077]  = 1;
  ram[11078]  = 1;
  ram[11079]  = 1;
  ram[11080]  = 1;
  ram[11081]  = 0;
  ram[11082]  = 0;
  ram[11083]  = 1;
  ram[11084]  = 1;
  ram[11085]  = 1;
  ram[11086]  = 1;
  ram[11087]  = 1;
  ram[11088]  = 1;
  ram[11089]  = 0;
  ram[11090]  = 0;
  ram[11091]  = 1;
  ram[11092]  = 1;
  ram[11093]  = 1;
  ram[11094]  = 1;
  ram[11095]  = 1;
  ram[11096]  = 1;
  ram[11097]  = 1;
  ram[11098]  = 1;
  ram[11099]  = 1;
  ram[11100]  = 1;
  ram[11101]  = 1;
  ram[11102]  = 1;
  ram[11103]  = 1;
  ram[11104]  = 1;
  ram[11105]  = 1;
  ram[11106]  = 1;
  ram[11107]  = 1;
  ram[11108]  = 1;
  ram[11109]  = 1;
  ram[11110]  = 1;
  ram[11111]  = 1;
  ram[11112]  = 1;
  ram[11113]  = 1;
  ram[11114]  = 1;
  ram[11115]  = 1;
  ram[11116]  = 1;
  ram[11117]  = 1;
  ram[11118]  = 0;
  ram[11119]  = 0;
  ram[11120]  = 0;
  ram[11121]  = 0;
  ram[11122]  = 0;
  ram[11123]  = 0;
  ram[11124]  = 0;
  ram[11125]  = 0;
  ram[11126]  = 1;
  ram[11127]  = 1;
  ram[11128]  = 0;
  ram[11129]  = 0;
  ram[11130]  = 0;
  ram[11131]  = 0;
  ram[11132]  = 0;
  ram[11133]  = 0;
  ram[11134]  = 0;
  ram[11135]  = 0;
  ram[11136]  = 0;
  ram[11137]  = 1;
  ram[11138]  = 1;
  ram[11139]  = 1;
  ram[11140]  = 1;
  ram[11141]  = 0;
  ram[11142]  = 1;
  ram[11143]  = 1;
  ram[11144]  = 1;
  ram[11145]  = 1;
  ram[11146]  = 0;
  ram[11147]  = 0;
  ram[11148]  = 1;
  ram[11149]  = 1;
  ram[11150]  = 1;
  ram[11151]  = 1;
  ram[11152]  = 1;
  ram[11153]  = 1;
  ram[11154]  = 1;
  ram[11155]  = 1;
  ram[11156]  = 1;
  ram[11157]  = 1;
  ram[11158]  = 1;
  ram[11159]  = 1;
  ram[11160]  = 1;
  ram[11161]  = 1;
  ram[11162]  = 1;
  ram[11163]  = 1;
  ram[11164]  = 1;
  ram[11165]  = 1;
  ram[11166]  = 1;
  ram[11167]  = 1;
  ram[11168]  = 1;
  ram[11169]  = 0;
  ram[11170]  = 0;
  ram[11171]  = 1;
  ram[11172]  = 1;
  ram[11173]  = 1;
  ram[11174]  = 1;
  ram[11175]  = 1;
  ram[11176]  = 1;
  ram[11177]  = 1;
  ram[11178]  = 1;
  ram[11179]  = 1;
  ram[11180]  = 1;
  ram[11181]  = 1;
  ram[11182]  = 1;
  ram[11183]  = 1;
  ram[11184]  = 1;
  ram[11185]  = 1;
  ram[11186]  = 1;
  ram[11187]  = 1;
  ram[11188]  = 1;
  ram[11189]  = 1;
  ram[11190]  = 1;
  ram[11191]  = 1;
  ram[11192]  = 1;
  ram[11193]  = 1;
  ram[11194]  = 1;
  ram[11195]  = 1;
  ram[11196]  = 1;
  ram[11197]  = 1;
  ram[11198]  = 1;
  ram[11199]  = 1;
  ram[11200]  = 1;
  ram[11201]  = 1;
  ram[11202]  = 1;
  ram[11203]  = 1;
  ram[11204]  = 1;
  ram[11205]  = 1;
  ram[11206]  = 1;
  ram[11207]  = 1;
  ram[11208]  = 1;
  ram[11209]  = 1;
  ram[11210]  = 1;
  ram[11211]  = 1;
  ram[11212]  = 1;
  ram[11213]  = 1;
  ram[11214]  = 1;
  ram[11215]  = 1;
  ram[11216]  = 1;
  ram[11217]  = 1;
  ram[11218]  = 1;
  ram[11219]  = 1;
  ram[11220]  = 0;
  ram[11221]  = 0;
  ram[11222]  = 0;
  ram[11223]  = 0;
  ram[11224]  = 0;
  ram[11225]  = 0;
  ram[11226]  = 0;
  ram[11227]  = 0;
  ram[11228]  = 1;
  ram[11229]  = 1;
  ram[11230]  = 1;
  ram[11231]  = 1;
  ram[11232]  = 1;
  ram[11233]  = 1;
  ram[11234]  = 1;
  ram[11235]  = 0;
  ram[11236]  = 1;
  ram[11237]  = 1;
  ram[11238]  = 1;
  ram[11239]  = 1;
  ram[11240]  = 1;
  ram[11241]  = 1;
  ram[11242]  = 0;
  ram[11243]  = 0;
  ram[11244]  = 0;
  ram[11245]  = 0;
  ram[11246]  = 0;
  ram[11247]  = 1;
  ram[11248]  = 1;
  ram[11249]  = 1;
  ram[11250]  = 1;
  ram[11251]  = 1;
  ram[11252]  = 0;
  ram[11253]  = 0;
  ram[11254]  = 1;
  ram[11255]  = 1;
  ram[11256]  = 1;
  ram[11257]  = 0;
  ram[11258]  = 0;
  ram[11259]  = 0;
  ram[11260]  = 0;
  ram[11261]  = 0;
  ram[11262]  = 0;
  ram[11263]  = 0;
  ram[11264]  = 0;
  ram[11265]  = 0;
  ram[11266]  = 1;
  ram[11267]  = 1;
  ram[11268]  = 1;
  ram[11269]  = 1;
  ram[11270]  = 1;
  ram[11271]  = 1;
  ram[11272]  = 0;
  ram[11273]  = 0;
  ram[11274]  = 1;
  ram[11275]  = 1;
  ram[11276]  = 1;
  ram[11277]  = 1;
  ram[11278]  = 1;
  ram[11279]  = 1;
  ram[11280]  = 1;
  ram[11281]  = 0;
  ram[11282]  = 0;
  ram[11283]  = 1;
  ram[11284]  = 1;
  ram[11285]  = 1;
  ram[11286]  = 1;
  ram[11287]  = 1;
  ram[11288]  = 0;
  ram[11289]  = 0;
  ram[11290]  = 1;
  ram[11291]  = 1;
  ram[11292]  = 1;
  ram[11293]  = 1;
  ram[11294]  = 1;
  ram[11295]  = 1;
  ram[11296]  = 1;
  ram[11297]  = 1;
  ram[11298]  = 1;
  ram[11299]  = 1;
  ram[11300]  = 1;
  ram[11301]  = 1;
  ram[11302]  = 1;
  ram[11303]  = 1;
  ram[11304]  = 1;
  ram[11305]  = 1;
  ram[11306]  = 1;
  ram[11307]  = 1;
  ram[11308]  = 1;
  ram[11309]  = 1;
  ram[11310]  = 1;
  ram[11311]  = 1;
  ram[11312]  = 1;
  ram[11313]  = 1;
  ram[11314]  = 1;
  ram[11315]  = 0;
  ram[11316]  = 0;
  ram[11317]  = 0;
  ram[11318]  = 0;
  ram[11319]  = 0;
  ram[11320]  = 0;
  ram[11321]  = 0;
  ram[11322]  = 0;
  ram[11323]  = 0;
  ram[11324]  = 1;
  ram[11325]  = 1;
  ram[11326]  = 1;
  ram[11327]  = 1;
  ram[11328]  = 0;
  ram[11329]  = 0;
  ram[11330]  = 1;
  ram[11331]  = 1;
  ram[11332]  = 1;
  ram[11333]  = 1;
  ram[11334]  = 1;
  ram[11335]  = 0;
  ram[11336]  = 0;
  ram[11337]  = 1;
  ram[11338]  = 1;
  ram[11339]  = 1;
  ram[11340]  = 1;
  ram[11341]  = 0;
  ram[11342]  = 1;
  ram[11343]  = 1;
  ram[11344]  = 1;
  ram[11345]  = 1;
  ram[11346]  = 0;
  ram[11347]  = 0;
  ram[11348]  = 1;
  ram[11349]  = 1;
  ram[11350]  = 1;
  ram[11351]  = 1;
  ram[11352]  = 1;
  ram[11353]  = 1;
  ram[11354]  = 1;
  ram[11355]  = 1;
  ram[11356]  = 1;
  ram[11357]  = 1;
  ram[11358]  = 1;
  ram[11359]  = 1;
  ram[11360]  = 1;
  ram[11361]  = 1;
  ram[11362]  = 1;
  ram[11363]  = 1;
  ram[11364]  = 1;
  ram[11365]  = 1;
  ram[11366]  = 1;
  ram[11367]  = 1;
  ram[11368]  = 1;
  ram[11369]  = 0;
  ram[11370]  = 0;
  ram[11371]  = 1;
  ram[11372]  = 1;
  ram[11373]  = 1;
  ram[11374]  = 1;
  ram[11375]  = 1;
  ram[11376]  = 1;
  ram[11377]  = 1;
  ram[11378]  = 1;
  ram[11379]  = 1;
  ram[11380]  = 1;
  ram[11381]  = 1;
  ram[11382]  = 1;
  ram[11383]  = 1;
  ram[11384]  = 1;
  ram[11385]  = 1;
  ram[11386]  = 1;
  ram[11387]  = 1;
  ram[11388]  = 1;
  ram[11389]  = 1;
  ram[11390]  = 1;
  ram[11391]  = 1;
  ram[11392]  = 1;
  ram[11393]  = 1;
  ram[11394]  = 1;
  ram[11395]  = 1;
  ram[11396]  = 1;
  ram[11397]  = 1;
  ram[11398]  = 1;
  ram[11399]  = 1;
  ram[11400]  = 1;
  ram[11401]  = 1;
  ram[11402]  = 1;
  ram[11403]  = 1;
  ram[11404]  = 1;
  ram[11405]  = 1;
  ram[11406]  = 1;
  ram[11407]  = 1;
  ram[11408]  = 1;
  ram[11409]  = 1;
  ram[11410]  = 1;
  ram[11411]  = 1;
  ram[11412]  = 1;
  ram[11413]  = 1;
  ram[11414]  = 1;
  ram[11415]  = 1;
  ram[11416]  = 1;
  ram[11417]  = 1;
  ram[11418]  = 1;
  ram[11419]  = 1;
  ram[11420]  = 0;
  ram[11421]  = 0;
  ram[11422]  = 1;
  ram[11423]  = 1;
  ram[11424]  = 1;
  ram[11425]  = 1;
  ram[11426]  = 1;
  ram[11427]  = 1;
  ram[11428]  = 1;
  ram[11429]  = 1;
  ram[11430]  = 1;
  ram[11431]  = 1;
  ram[11432]  = 1;
  ram[11433]  = 1;
  ram[11434]  = 1;
  ram[11435]  = 0;
  ram[11436]  = 1;
  ram[11437]  = 1;
  ram[11438]  = 1;
  ram[11439]  = 1;
  ram[11440]  = 1;
  ram[11441]  = 0;
  ram[11442]  = 0;
  ram[11443]  = 0;
  ram[11444]  = 0;
  ram[11445]  = 0;
  ram[11446]  = 0;
  ram[11447]  = 1;
  ram[11448]  = 1;
  ram[11449]  = 1;
  ram[11450]  = 1;
  ram[11451]  = 1;
  ram[11452]  = 0;
  ram[11453]  = 0;
  ram[11454]  = 1;
  ram[11455]  = 1;
  ram[11456]  = 1;
  ram[11457]  = 0;
  ram[11458]  = 0;
  ram[11459]  = 1;
  ram[11460]  = 1;
  ram[11461]  = 1;
  ram[11462]  = 1;
  ram[11463]  = 1;
  ram[11464]  = 1;
  ram[11465]  = 1;
  ram[11466]  = 1;
  ram[11467]  = 1;
  ram[11468]  = 1;
  ram[11469]  = 1;
  ram[11470]  = 1;
  ram[11471]  = 1;
  ram[11472]  = 0;
  ram[11473]  = 0;
  ram[11474]  = 1;
  ram[11475]  = 1;
  ram[11476]  = 1;
  ram[11477]  = 1;
  ram[11478]  = 1;
  ram[11479]  = 1;
  ram[11480]  = 1;
  ram[11481]  = 0;
  ram[11482]  = 0;
  ram[11483]  = 1;
  ram[11484]  = 1;
  ram[11485]  = 1;
  ram[11486]  = 1;
  ram[11487]  = 1;
  ram[11488]  = 0;
  ram[11489]  = 0;
  ram[11490]  = 1;
  ram[11491]  = 1;
  ram[11492]  = 1;
  ram[11493]  = 1;
  ram[11494]  = 1;
  ram[11495]  = 1;
  ram[11496]  = 1;
  ram[11497]  = 1;
  ram[11498]  = 1;
  ram[11499]  = 1;
  ram[11500]  = 1;
  ram[11501]  = 1;
  ram[11502]  = 1;
  ram[11503]  = 1;
  ram[11504]  = 1;
  ram[11505]  = 1;
  ram[11506]  = 1;
  ram[11507]  = 1;
  ram[11508]  = 1;
  ram[11509]  = 1;
  ram[11510]  = 1;
  ram[11511]  = 1;
  ram[11512]  = 1;
  ram[11513]  = 1;
  ram[11514]  = 1;
  ram[11515]  = 0;
  ram[11516]  = 0;
  ram[11517]  = 1;
  ram[11518]  = 1;
  ram[11519]  = 1;
  ram[11520]  = 1;
  ram[11521]  = 0;
  ram[11522]  = 0;
  ram[11523]  = 1;
  ram[11524]  = 1;
  ram[11525]  = 1;
  ram[11526]  = 1;
  ram[11527]  = 1;
  ram[11528]  = 0;
  ram[11529]  = 0;
  ram[11530]  = 1;
  ram[11531]  = 1;
  ram[11532]  = 1;
  ram[11533]  = 1;
  ram[11534]  = 1;
  ram[11535]  = 0;
  ram[11536]  = 0;
  ram[11537]  = 1;
  ram[11538]  = 1;
  ram[11539]  = 1;
  ram[11540]  = 1;
  ram[11541]  = 1;
  ram[11542]  = 1;
  ram[11543]  = 1;
  ram[11544]  = 1;
  ram[11545]  = 1;
  ram[11546]  = 0;
  ram[11547]  = 0;
  ram[11548]  = 1;
  ram[11549]  = 1;
  ram[11550]  = 1;
  ram[11551]  = 1;
  ram[11552]  = 1;
  ram[11553]  = 1;
  ram[11554]  = 1;
  ram[11555]  = 1;
  ram[11556]  = 1;
  ram[11557]  = 1;
  ram[11558]  = 1;
  ram[11559]  = 1;
  ram[11560]  = 1;
  ram[11561]  = 1;
  ram[11562]  = 1;
  ram[11563]  = 1;
  ram[11564]  = 1;
  ram[11565]  = 1;
  ram[11566]  = 1;
  ram[11567]  = 1;
  ram[11568]  = 1;
  ram[11569]  = 0;
  ram[11570]  = 0;
  ram[11571]  = 1;
  ram[11572]  = 1;
  ram[11573]  = 1;
  ram[11574]  = 1;
  ram[11575]  = 1;
  ram[11576]  = 1;
  ram[11577]  = 1;
  ram[11578]  = 1;
  ram[11579]  = 1;
  ram[11580]  = 1;
  ram[11581]  = 1;
  ram[11582]  = 1;
  ram[11583]  = 1;
  ram[11584]  = 1;
  ram[11585]  = 1;
  ram[11586]  = 1;
  ram[11587]  = 1;
  ram[11588]  = 1;
  ram[11589]  = 1;
  ram[11590]  = 1;
  ram[11591]  = 1;
  ram[11592]  = 1;
  ram[11593]  = 1;
  ram[11594]  = 1;
  ram[11595]  = 1;
  ram[11596]  = 1;
  ram[11597]  = 1;
  ram[11598]  = 1;
  ram[11599]  = 1;
  ram[11600]  = 1;
  ram[11601]  = 1;
  ram[11602]  = 1;
  ram[11603]  = 1;
  ram[11604]  = 1;
  ram[11605]  = 1;
  ram[11606]  = 1;
  ram[11607]  = 1;
  ram[11608]  = 1;
  ram[11609]  = 1;
  ram[11610]  = 1;
  ram[11611]  = 1;
  ram[11612]  = 1;
  ram[11613]  = 1;
  ram[11614]  = 1;
  ram[11615]  = 1;
  ram[11616]  = 1;
  ram[11617]  = 1;
  ram[11618]  = 1;
  ram[11619]  = 1;
  ram[11620]  = 0;
  ram[11621]  = 0;
  ram[11622]  = 1;
  ram[11623]  = 1;
  ram[11624]  = 1;
  ram[11625]  = 1;
  ram[11626]  = 1;
  ram[11627]  = 1;
  ram[11628]  = 1;
  ram[11629]  = 1;
  ram[11630]  = 1;
  ram[11631]  = 1;
  ram[11632]  = 1;
  ram[11633]  = 1;
  ram[11634]  = 1;
  ram[11635]  = 0;
  ram[11636]  = 1;
  ram[11637]  = 1;
  ram[11638]  = 1;
  ram[11639]  = 1;
  ram[11640]  = 0;
  ram[11641]  = 0;
  ram[11642]  = 0;
  ram[11643]  = 1;
  ram[11644]  = 1;
  ram[11645]  = 0;
  ram[11646]  = 0;
  ram[11647]  = 1;
  ram[11648]  = 1;
  ram[11649]  = 1;
  ram[11650]  = 1;
  ram[11651]  = 1;
  ram[11652]  = 0;
  ram[11653]  = 0;
  ram[11654]  = 1;
  ram[11655]  = 1;
  ram[11656]  = 1;
  ram[11657]  = 0;
  ram[11658]  = 0;
  ram[11659]  = 1;
  ram[11660]  = 1;
  ram[11661]  = 1;
  ram[11662]  = 1;
  ram[11663]  = 1;
  ram[11664]  = 1;
  ram[11665]  = 1;
  ram[11666]  = 1;
  ram[11667]  = 1;
  ram[11668]  = 1;
  ram[11669]  = 1;
  ram[11670]  = 1;
  ram[11671]  = 1;
  ram[11672]  = 0;
  ram[11673]  = 0;
  ram[11674]  = 1;
  ram[11675]  = 1;
  ram[11676]  = 1;
  ram[11677]  = 1;
  ram[11678]  = 1;
  ram[11679]  = 1;
  ram[11680]  = 1;
  ram[11681]  = 0;
  ram[11682]  = 0;
  ram[11683]  = 1;
  ram[11684]  = 1;
  ram[11685]  = 1;
  ram[11686]  = 1;
  ram[11687]  = 1;
  ram[11688]  = 0;
  ram[11689]  = 0;
  ram[11690]  = 1;
  ram[11691]  = 1;
  ram[11692]  = 1;
  ram[11693]  = 1;
  ram[11694]  = 1;
  ram[11695]  = 1;
  ram[11696]  = 1;
  ram[11697]  = 1;
  ram[11698]  = 1;
  ram[11699]  = 1;
  ram[11700]  = 1;
  ram[11701]  = 1;
  ram[11702]  = 1;
  ram[11703]  = 1;
  ram[11704]  = 1;
  ram[11705]  = 1;
  ram[11706]  = 1;
  ram[11707]  = 1;
  ram[11708]  = 1;
  ram[11709]  = 1;
  ram[11710]  = 1;
  ram[11711]  = 1;
  ram[11712]  = 1;
  ram[11713]  = 1;
  ram[11714]  = 1;
  ram[11715]  = 1;
  ram[11716]  = 1;
  ram[11717]  = 1;
  ram[11718]  = 1;
  ram[11719]  = 1;
  ram[11720]  = 1;
  ram[11721]  = 0;
  ram[11722]  = 0;
  ram[11723]  = 1;
  ram[11724]  = 1;
  ram[11725]  = 1;
  ram[11726]  = 1;
  ram[11727]  = 1;
  ram[11728]  = 0;
  ram[11729]  = 0;
  ram[11730]  = 1;
  ram[11731]  = 1;
  ram[11732]  = 1;
  ram[11733]  = 1;
  ram[11734]  = 1;
  ram[11735]  = 0;
  ram[11736]  = 0;
  ram[11737]  = 1;
  ram[11738]  = 1;
  ram[11739]  = 1;
  ram[11740]  = 1;
  ram[11741]  = 1;
  ram[11742]  = 1;
  ram[11743]  = 1;
  ram[11744]  = 1;
  ram[11745]  = 1;
  ram[11746]  = 0;
  ram[11747]  = 0;
  ram[11748]  = 1;
  ram[11749]  = 1;
  ram[11750]  = 1;
  ram[11751]  = 1;
  ram[11752]  = 1;
  ram[11753]  = 1;
  ram[11754]  = 1;
  ram[11755]  = 1;
  ram[11756]  = 1;
  ram[11757]  = 1;
  ram[11758]  = 1;
  ram[11759]  = 1;
  ram[11760]  = 1;
  ram[11761]  = 1;
  ram[11762]  = 1;
  ram[11763]  = 1;
  ram[11764]  = 1;
  ram[11765]  = 1;
  ram[11766]  = 1;
  ram[11767]  = 1;
  ram[11768]  = 1;
  ram[11769]  = 0;
  ram[11770]  = 0;
  ram[11771]  = 1;
  ram[11772]  = 1;
  ram[11773]  = 1;
  ram[11774]  = 1;
  ram[11775]  = 1;
  ram[11776]  = 1;
  ram[11777]  = 1;
  ram[11778]  = 1;
  ram[11779]  = 1;
  ram[11780]  = 1;
  ram[11781]  = 1;
  ram[11782]  = 1;
  ram[11783]  = 1;
  ram[11784]  = 1;
  ram[11785]  = 1;
  ram[11786]  = 1;
  ram[11787]  = 1;
  ram[11788]  = 1;
  ram[11789]  = 1;
  ram[11790]  = 1;
  ram[11791]  = 1;
  ram[11792]  = 1;
  ram[11793]  = 1;
  ram[11794]  = 1;
  ram[11795]  = 1;
  ram[11796]  = 1;
  ram[11797]  = 1;
  ram[11798]  = 1;
  ram[11799]  = 1;
  ram[11800]  = 1;
  ram[11801]  = 1;
  ram[11802]  = 1;
  ram[11803]  = 1;
  ram[11804]  = 1;
  ram[11805]  = 1;
  ram[11806]  = 1;
  ram[11807]  = 1;
  ram[11808]  = 1;
  ram[11809]  = 1;
  ram[11810]  = 1;
  ram[11811]  = 1;
  ram[11812]  = 1;
  ram[11813]  = 1;
  ram[11814]  = 1;
  ram[11815]  = 1;
  ram[11816]  = 1;
  ram[11817]  = 1;
  ram[11818]  = 1;
  ram[11819]  = 1;
  ram[11820]  = 0;
  ram[11821]  = 0;
  ram[11822]  = 1;
  ram[11823]  = 1;
  ram[11824]  = 1;
  ram[11825]  = 1;
  ram[11826]  = 1;
  ram[11827]  = 1;
  ram[11828]  = 1;
  ram[11829]  = 1;
  ram[11830]  = 1;
  ram[11831]  = 1;
  ram[11832]  = 1;
  ram[11833]  = 1;
  ram[11834]  = 1;
  ram[11835]  = 0;
  ram[11836]  = 1;
  ram[11837]  = 1;
  ram[11838]  = 0;
  ram[11839]  = 0;
  ram[11840]  = 0;
  ram[11841]  = 0;
  ram[11842]  = 1;
  ram[11843]  = 1;
  ram[11844]  = 1;
  ram[11845]  = 1;
  ram[11846]  = 0;
  ram[11847]  = 0;
  ram[11848]  = 1;
  ram[11849]  = 1;
  ram[11850]  = 1;
  ram[11851]  = 1;
  ram[11852]  = 0;
  ram[11853]  = 0;
  ram[11854]  = 1;
  ram[11855]  = 1;
  ram[11856]  = 1;
  ram[11857]  = 0;
  ram[11858]  = 0;
  ram[11859]  = 1;
  ram[11860]  = 1;
  ram[11861]  = 1;
  ram[11862]  = 1;
  ram[11863]  = 1;
  ram[11864]  = 1;
  ram[11865]  = 1;
  ram[11866]  = 1;
  ram[11867]  = 1;
  ram[11868]  = 1;
  ram[11869]  = 1;
  ram[11870]  = 1;
  ram[11871]  = 1;
  ram[11872]  = 0;
  ram[11873]  = 0;
  ram[11874]  = 1;
  ram[11875]  = 1;
  ram[11876]  = 1;
  ram[11877]  = 1;
  ram[11878]  = 1;
  ram[11879]  = 1;
  ram[11880]  = 1;
  ram[11881]  = 0;
  ram[11882]  = 0;
  ram[11883]  = 1;
  ram[11884]  = 1;
  ram[11885]  = 1;
  ram[11886]  = 1;
  ram[11887]  = 1;
  ram[11888]  = 0;
  ram[11889]  = 0;
  ram[11890]  = 1;
  ram[11891]  = 1;
  ram[11892]  = 1;
  ram[11893]  = 1;
  ram[11894]  = 1;
  ram[11895]  = 1;
  ram[11896]  = 1;
  ram[11897]  = 1;
  ram[11898]  = 1;
  ram[11899]  = 1;
  ram[11900]  = 1;
  ram[11901]  = 1;
  ram[11902]  = 1;
  ram[11903]  = 1;
  ram[11904]  = 1;
  ram[11905]  = 1;
  ram[11906]  = 1;
  ram[11907]  = 1;
  ram[11908]  = 1;
  ram[11909]  = 1;
  ram[11910]  = 1;
  ram[11911]  = 1;
  ram[11912]  = 1;
  ram[11913]  = 1;
  ram[11914]  = 1;
  ram[11915]  = 1;
  ram[11916]  = 1;
  ram[11917]  = 1;
  ram[11918]  = 1;
  ram[11919]  = 1;
  ram[11920]  = 1;
  ram[11921]  = 0;
  ram[11922]  = 0;
  ram[11923]  = 1;
  ram[11924]  = 1;
  ram[11925]  = 1;
  ram[11926]  = 1;
  ram[11927]  = 1;
  ram[11928]  = 0;
  ram[11929]  = 0;
  ram[11930]  = 1;
  ram[11931]  = 1;
  ram[11932]  = 1;
  ram[11933]  = 1;
  ram[11934]  = 1;
  ram[11935]  = 0;
  ram[11936]  = 0;
  ram[11937]  = 1;
  ram[11938]  = 1;
  ram[11939]  = 1;
  ram[11940]  = 1;
  ram[11941]  = 1;
  ram[11942]  = 1;
  ram[11943]  = 1;
  ram[11944]  = 1;
  ram[11945]  = 1;
  ram[11946]  = 0;
  ram[11947]  = 0;
  ram[11948]  = 1;
  ram[11949]  = 1;
  ram[11950]  = 1;
  ram[11951]  = 1;
  ram[11952]  = 1;
  ram[11953]  = 1;
  ram[11954]  = 1;
  ram[11955]  = 1;
  ram[11956]  = 1;
  ram[11957]  = 1;
  ram[11958]  = 1;
  ram[11959]  = 1;
  ram[11960]  = 1;
  ram[11961]  = 1;
  ram[11962]  = 1;
  ram[11963]  = 1;
  ram[11964]  = 1;
  ram[11965]  = 1;
  ram[11966]  = 1;
  ram[11967]  = 1;
  ram[11968]  = 0;
  ram[11969]  = 0;
  ram[11970]  = 0;
  ram[11971]  = 1;
  ram[11972]  = 1;
  ram[11973]  = 1;
  ram[11974]  = 1;
  ram[11975]  = 1;
  ram[11976]  = 1;
  ram[11977]  = 1;
  ram[11978]  = 1;
  ram[11979]  = 1;
  ram[11980]  = 1;
  ram[11981]  = 1;
  ram[11982]  = 1;
  ram[11983]  = 1;
  ram[11984]  = 1;
  ram[11985]  = 1;
  ram[11986]  = 1;
  ram[11987]  = 1;
  ram[11988]  = 1;
  ram[11989]  = 1;
  ram[11990]  = 1;
  ram[11991]  = 1;
  ram[11992]  = 1;
  ram[11993]  = 1;
  ram[11994]  = 1;
  ram[11995]  = 1;
  ram[11996]  = 1;
  ram[11997]  = 1;
  ram[11998]  = 1;
  ram[11999]  = 1;
  ram[12000]  = 1;
  ram[12001]  = 1;
  ram[12002]  = 1;
  ram[12003]  = 1;
  ram[12004]  = 1;
  ram[12005]  = 1;
  ram[12006]  = 1;
  ram[12007]  = 1;
  ram[12008]  = 1;
  ram[12009]  = 1;
  ram[12010]  = 1;
  ram[12011]  = 1;
  ram[12012]  = 1;
  ram[12013]  = 1;
  ram[12014]  = 1;
  ram[12015]  = 1;
  ram[12016]  = 1;
  ram[12017]  = 1;
  ram[12018]  = 1;
  ram[12019]  = 1;
  ram[12020]  = 1;
  ram[12021]  = 1;
  ram[12022]  = 1;
  ram[12023]  = 1;
  ram[12024]  = 1;
  ram[12025]  = 1;
  ram[12026]  = 1;
  ram[12027]  = 1;
  ram[12028]  = 1;
  ram[12029]  = 1;
  ram[12030]  = 1;
  ram[12031]  = 1;
  ram[12032]  = 1;
  ram[12033]  = 1;
  ram[12034]  = 1;
  ram[12035]  = 0;
  ram[12036]  = 1;
  ram[12037]  = 1;
  ram[12038]  = 1;
  ram[12039]  = 0;
  ram[12040]  = 1;
  ram[12041]  = 1;
  ram[12042]  = 1;
  ram[12043]  = 1;
  ram[12044]  = 1;
  ram[12045]  = 1;
  ram[12046]  = 0;
  ram[12047]  = 0;
  ram[12048]  = 1;
  ram[12049]  = 1;
  ram[12050]  = 1;
  ram[12051]  = 1;
  ram[12052]  = 0;
  ram[12053]  = 0;
  ram[12054]  = 1;
  ram[12055]  = 1;
  ram[12056]  = 1;
  ram[12057]  = 1;
  ram[12058]  = 1;
  ram[12059]  = 1;
  ram[12060]  = 1;
  ram[12061]  = 1;
  ram[12062]  = 1;
  ram[12063]  = 1;
  ram[12064]  = 1;
  ram[12065]  = 1;
  ram[12066]  = 1;
  ram[12067]  = 1;
  ram[12068]  = 1;
  ram[12069]  = 1;
  ram[12070]  = 1;
  ram[12071]  = 1;
  ram[12072]  = 0;
  ram[12073]  = 0;
  ram[12074]  = 1;
  ram[12075]  = 1;
  ram[12076]  = 1;
  ram[12077]  = 1;
  ram[12078]  = 1;
  ram[12079]  = 1;
  ram[12080]  = 1;
  ram[12081]  = 0;
  ram[12082]  = 0;
  ram[12083]  = 1;
  ram[12084]  = 1;
  ram[12085]  = 1;
  ram[12086]  = 1;
  ram[12087]  = 1;
  ram[12088]  = 0;
  ram[12089]  = 0;
  ram[12090]  = 1;
  ram[12091]  = 1;
  ram[12092]  = 1;
  ram[12093]  = 1;
  ram[12094]  = 1;
  ram[12095]  = 1;
  ram[12096]  = 1;
  ram[12097]  = 1;
  ram[12098]  = 1;
  ram[12099]  = 1;
  ram[12100]  = 1;
  ram[12101]  = 1;
  ram[12102]  = 1;
  ram[12103]  = 1;
  ram[12104]  = 1;
  ram[12105]  = 1;
  ram[12106]  = 1;
  ram[12107]  = 1;
  ram[12108]  = 1;
  ram[12109]  = 1;
  ram[12110]  = 1;
  ram[12111]  = 1;
  ram[12112]  = 1;
  ram[12113]  = 1;
  ram[12114]  = 1;
  ram[12115]  = 1;
  ram[12116]  = 1;
  ram[12117]  = 1;
  ram[12118]  = 1;
  ram[12119]  = 1;
  ram[12120]  = 1;
  ram[12121]  = 0;
  ram[12122]  = 0;
  ram[12123]  = 1;
  ram[12124]  = 1;
  ram[12125]  = 1;
  ram[12126]  = 1;
  ram[12127]  = 1;
  ram[12128]  = 0;
  ram[12129]  = 0;
  ram[12130]  = 1;
  ram[12131]  = 1;
  ram[12132]  = 1;
  ram[12133]  = 1;
  ram[12134]  = 1;
  ram[12135]  = 0;
  ram[12136]  = 0;
  ram[12137]  = 1;
  ram[12138]  = 1;
  ram[12139]  = 1;
  ram[12140]  = 1;
  ram[12141]  = 1;
  ram[12142]  = 1;
  ram[12143]  = 1;
  ram[12144]  = 1;
  ram[12145]  = 1;
  ram[12146]  = 0;
  ram[12147]  = 0;
  ram[12148]  = 1;
  ram[12149]  = 1;
  ram[12150]  = 1;
  ram[12151]  = 1;
  ram[12152]  = 1;
  ram[12153]  = 1;
  ram[12154]  = 1;
  ram[12155]  = 1;
  ram[12156]  = 1;
  ram[12157]  = 1;
  ram[12158]  = 1;
  ram[12159]  = 1;
  ram[12160]  = 1;
  ram[12161]  = 1;
  ram[12162]  = 1;
  ram[12163]  = 1;
  ram[12164]  = 1;
  ram[12165]  = 1;
  ram[12166]  = 1;
  ram[12167]  = 0;
  ram[12168]  = 0;
  ram[12169]  = 0;
  ram[12170]  = 0;
  ram[12171]  = 1;
  ram[12172]  = 1;
  ram[12173]  = 1;
  ram[12174]  = 1;
  ram[12175]  = 1;
  ram[12176]  = 1;
  ram[12177]  = 1;
  ram[12178]  = 1;
  ram[12179]  = 1;
  ram[12180]  = 1;
  ram[12181]  = 1;
  ram[12182]  = 1;
  ram[12183]  = 1;
  ram[12184]  = 1;
  ram[12185]  = 1;
  ram[12186]  = 1;
  ram[12187]  = 1;
  ram[12188]  = 1;
  ram[12189]  = 1;
  ram[12190]  = 1;
  ram[12191]  = 1;
  ram[12192]  = 1;
  ram[12193]  = 1;
  ram[12194]  = 1;
  ram[12195]  = 1;
  ram[12196]  = 1;
  ram[12197]  = 1;
  ram[12198]  = 1;
  ram[12199]  = 1;
  ram[12200]  = 1;
  ram[12201]  = 1;
  ram[12202]  = 1;
  ram[12203]  = 1;
  ram[12204]  = 1;
  ram[12205]  = 1;
  ram[12206]  = 1;
  ram[12207]  = 1;
  ram[12208]  = 1;
  ram[12209]  = 1;
  ram[12210]  = 1;
  ram[12211]  = 1;
  ram[12212]  = 1;
  ram[12213]  = 1;
  ram[12214]  = 1;
  ram[12215]  = 1;
  ram[12216]  = 1;
  ram[12217]  = 1;
  ram[12218]  = 1;
  ram[12219]  = 1;
  ram[12220]  = 1;
  ram[12221]  = 1;
  ram[12222]  = 1;
  ram[12223]  = 1;
  ram[12224]  = 1;
  ram[12225]  = 1;
  ram[12226]  = 1;
  ram[12227]  = 1;
  ram[12228]  = 1;
  ram[12229]  = 1;
  ram[12230]  = 1;
  ram[12231]  = 1;
  ram[12232]  = 1;
  ram[12233]  = 1;
  ram[12234]  = 0;
  ram[12235]  = 0;
  ram[12236]  = 1;
  ram[12237]  = 1;
  ram[12238]  = 1;
  ram[12239]  = 1;
  ram[12240]  = 1;
  ram[12241]  = 1;
  ram[12242]  = 1;
  ram[12243]  = 1;
  ram[12244]  = 1;
  ram[12245]  = 1;
  ram[12246]  = 1;
  ram[12247]  = 0;
  ram[12248]  = 0;
  ram[12249]  = 1;
  ram[12250]  = 1;
  ram[12251]  = 0;
  ram[12252]  = 0;
  ram[12253]  = 1;
  ram[12254]  = 1;
  ram[12255]  = 1;
  ram[12256]  = 1;
  ram[12257]  = 1;
  ram[12258]  = 1;
  ram[12259]  = 1;
  ram[12260]  = 1;
  ram[12261]  = 1;
  ram[12262]  = 1;
  ram[12263]  = 1;
  ram[12264]  = 1;
  ram[12265]  = 1;
  ram[12266]  = 1;
  ram[12267]  = 0;
  ram[12268]  = 1;
  ram[12269]  = 1;
  ram[12270]  = 1;
  ram[12271]  = 0;
  ram[12272]  = 0;
  ram[12273]  = 0;
  ram[12274]  = 1;
  ram[12275]  = 1;
  ram[12276]  = 1;
  ram[12277]  = 1;
  ram[12278]  = 1;
  ram[12279]  = 1;
  ram[12280]  = 1;
  ram[12281]  = 1;
  ram[12282]  = 0;
  ram[12283]  = 0;
  ram[12284]  = 0;
  ram[12285]  = 0;
  ram[12286]  = 0;
  ram[12287]  = 0;
  ram[12288]  = 0;
  ram[12289]  = 0;
  ram[12290]  = 1;
  ram[12291]  = 1;
  ram[12292]  = 1;
  ram[12293]  = 1;
  ram[12294]  = 1;
  ram[12295]  = 1;
  ram[12296]  = 1;
  ram[12297]  = 1;
  ram[12298]  = 1;
  ram[12299]  = 1;
  ram[12300]  = 1;
  ram[12301]  = 1;
  ram[12302]  = 1;
  ram[12303]  = 1;
  ram[12304]  = 1;
  ram[12305]  = 1;
  ram[12306]  = 1;
  ram[12307]  = 1;
  ram[12308]  = 1;
  ram[12309]  = 1;
  ram[12310]  = 1;
  ram[12311]  = 1;
  ram[12312]  = 1;
  ram[12313]  = 1;
  ram[12314]  = 1;
  ram[12315]  = 1;
  ram[12316]  = 1;
  ram[12317]  = 1;
  ram[12318]  = 1;
  ram[12319]  = 1;
  ram[12320]  = 1;
  ram[12321]  = 0;
  ram[12322]  = 0;
  ram[12323]  = 1;
  ram[12324]  = 1;
  ram[12325]  = 1;
  ram[12326]  = 1;
  ram[12327]  = 1;
  ram[12328]  = 0;
  ram[12329]  = 0;
  ram[12330]  = 1;
  ram[12331]  = 1;
  ram[12332]  = 1;
  ram[12333]  = 1;
  ram[12334]  = 1;
  ram[12335]  = 0;
  ram[12336]  = 0;
  ram[12337]  = 1;
  ram[12338]  = 1;
  ram[12339]  = 1;
  ram[12340]  = 1;
  ram[12341]  = 1;
  ram[12342]  = 1;
  ram[12343]  = 1;
  ram[12344]  = 1;
  ram[12345]  = 1;
  ram[12346]  = 0;
  ram[12347]  = 0;
  ram[12348]  = 1;
  ram[12349]  = 1;
  ram[12350]  = 1;
  ram[12351]  = 1;
  ram[12352]  = 1;
  ram[12353]  = 1;
  ram[12354]  = 1;
  ram[12355]  = 1;
  ram[12356]  = 1;
  ram[12357]  = 1;
  ram[12358]  = 1;
  ram[12359]  = 0;
  ram[12360]  = 0;
  ram[12361]  = 0;
  ram[12362]  = 0;
  ram[12363]  = 0;
  ram[12364]  = 0;
  ram[12365]  = 0;
  ram[12366]  = 0;
  ram[12367]  = 0;
  ram[12368]  = 0;
  ram[12369]  = 0;
  ram[12370]  = 1;
  ram[12371]  = 1;
  ram[12372]  = 1;
  ram[12373]  = 1;
  ram[12374]  = 1;
  ram[12375]  = 1;
  ram[12376]  = 1;
  ram[12377]  = 1;
  ram[12378]  = 1;
  ram[12379]  = 1;
  ram[12380]  = 1;
  ram[12381]  = 1;
  ram[12382]  = 1;
  ram[12383]  = 1;
  ram[12384]  = 1;
  ram[12385]  = 1;
  ram[12386]  = 1;
  ram[12387]  = 1;
  ram[12388]  = 1;
  ram[12389]  = 1;
  ram[12390]  = 1;
  ram[12391]  = 1;
  ram[12392]  = 1;
  ram[12393]  = 1;
  ram[12394]  = 1;
  ram[12395]  = 1;
  ram[12396]  = 1;
  ram[12397]  = 1;
  ram[12398]  = 1;
  ram[12399]  = 1;
  ram[12400]  = 1;
  ram[12401]  = 1;
  ram[12402]  = 1;
  ram[12403]  = 1;
  ram[12404]  = 1;
  ram[12405]  = 1;
  ram[12406]  = 1;
  ram[12407]  = 1;
  ram[12408]  = 1;
  ram[12409]  = 1;
  ram[12410]  = 1;
  ram[12411]  = 1;
  ram[12412]  = 1;
  ram[12413]  = 1;
  ram[12414]  = 1;
  ram[12415]  = 1;
  ram[12416]  = 1;
  ram[12417]  = 1;
  ram[12418]  = 1;
  ram[12419]  = 1;
  ram[12420]  = 1;
  ram[12421]  = 1;
  ram[12422]  = 1;
  ram[12423]  = 1;
  ram[12424]  = 1;
  ram[12425]  = 1;
  ram[12426]  = 1;
  ram[12427]  = 1;
  ram[12428]  = 1;
  ram[12429]  = 0;
  ram[12430]  = 0;
  ram[12431]  = 0;
  ram[12432]  = 0;
  ram[12433]  = 0;
  ram[12434]  = 0;
  ram[12435]  = 0;
  ram[12436]  = 1;
  ram[12437]  = 1;
  ram[12438]  = 1;
  ram[12439]  = 1;
  ram[12440]  = 1;
  ram[12441]  = 1;
  ram[12442]  = 1;
  ram[12443]  = 1;
  ram[12444]  = 1;
  ram[12445]  = 1;
  ram[12446]  = 1;
  ram[12447]  = 0;
  ram[12448]  = 0;
  ram[12449]  = 0;
  ram[12450]  = 0;
  ram[12451]  = 0;
  ram[12452]  = 0;
  ram[12453]  = 1;
  ram[12454]  = 1;
  ram[12455]  = 1;
  ram[12456]  = 1;
  ram[12457]  = 1;
  ram[12458]  = 1;
  ram[12459]  = 1;
  ram[12460]  = 1;
  ram[12461]  = 1;
  ram[12462]  = 1;
  ram[12463]  = 1;
  ram[12464]  = 1;
  ram[12465]  = 1;
  ram[12466]  = 1;
  ram[12467]  = 0;
  ram[12468]  = 0;
  ram[12469]  = 0;
  ram[12470]  = 0;
  ram[12471]  = 0;
  ram[12472]  = 0;
  ram[12473]  = 0;
  ram[12474]  = 1;
  ram[12475]  = 1;
  ram[12476]  = 1;
  ram[12477]  = 1;
  ram[12478]  = 1;
  ram[12479]  = 1;
  ram[12480]  = 1;
  ram[12481]  = 1;
  ram[12482]  = 0;
  ram[12483]  = 0;
  ram[12484]  = 0;
  ram[12485]  = 0;
  ram[12486]  = 0;
  ram[12487]  = 0;
  ram[12488]  = 0;
  ram[12489]  = 1;
  ram[12490]  = 1;
  ram[12491]  = 1;
  ram[12492]  = 1;
  ram[12493]  = 1;
  ram[12494]  = 1;
  ram[12495]  = 1;
  ram[12496]  = 1;
  ram[12497]  = 1;
  ram[12498]  = 1;
  ram[12499]  = 1;
  ram[12500]  = 1;
  ram[12501]  = 1;
  ram[12502]  = 1;
  ram[12503]  = 1;
  ram[12504]  = 1;
  ram[12505]  = 1;
  ram[12506]  = 1;
  ram[12507]  = 1;
  ram[12508]  = 1;
  ram[12509]  = 1;
  ram[12510]  = 1;
  ram[12511]  = 1;
  ram[12512]  = 1;
  ram[12513]  = 1;
  ram[12514]  = 1;
  ram[12515]  = 1;
  ram[12516]  = 1;
  ram[12517]  = 1;
  ram[12518]  = 1;
  ram[12519]  = 1;
  ram[12520]  = 1;
  ram[12521]  = 0;
  ram[12522]  = 0;
  ram[12523]  = 1;
  ram[12524]  = 1;
  ram[12525]  = 1;
  ram[12526]  = 1;
  ram[12527]  = 1;
  ram[12528]  = 0;
  ram[12529]  = 0;
  ram[12530]  = 1;
  ram[12531]  = 1;
  ram[12532]  = 1;
  ram[12533]  = 1;
  ram[12534]  = 1;
  ram[12535]  = 0;
  ram[12536]  = 0;
  ram[12537]  = 1;
  ram[12538]  = 1;
  ram[12539]  = 1;
  ram[12540]  = 1;
  ram[12541]  = 0;
  ram[12542]  = 0;
  ram[12543]  = 1;
  ram[12544]  = 0;
  ram[12545]  = 0;
  ram[12546]  = 0;
  ram[12547]  = 0;
  ram[12548]  = 1;
  ram[12549]  = 1;
  ram[12550]  = 1;
  ram[12551]  = 1;
  ram[12552]  = 1;
  ram[12553]  = 1;
  ram[12554]  = 1;
  ram[12555]  = 1;
  ram[12556]  = 1;
  ram[12557]  = 1;
  ram[12558]  = 1;
  ram[12559]  = 1;
  ram[12560]  = 0;
  ram[12561]  = 0;
  ram[12562]  = 0;
  ram[12563]  = 0;
  ram[12564]  = 0;
  ram[12565]  = 0;
  ram[12566]  = 0;
  ram[12567]  = 0;
  ram[12568]  = 0;
  ram[12569]  = 1;
  ram[12570]  = 1;
  ram[12571]  = 1;
  ram[12572]  = 1;
  ram[12573]  = 1;
  ram[12574]  = 1;
  ram[12575]  = 1;
  ram[12576]  = 1;
  ram[12577]  = 1;
  ram[12578]  = 1;
  ram[12579]  = 1;
  ram[12580]  = 1;
  ram[12581]  = 1;
  ram[12582]  = 1;
  ram[12583]  = 1;
  ram[12584]  = 1;
  ram[12585]  = 1;
  ram[12586]  = 1;
  ram[12587]  = 1;
  ram[12588]  = 1;
  ram[12589]  = 1;
  ram[12590]  = 1;
  ram[12591]  = 1;
  ram[12592]  = 1;
  ram[12593]  = 1;
  ram[12594]  = 1;
  ram[12595]  = 1;
  ram[12596]  = 1;
  ram[12597]  = 1;
  ram[12598]  = 1;
  ram[12599]  = 1;
  ram[12600]  = 1;
  ram[12601]  = 1;
  ram[12602]  = 1;
  ram[12603]  = 1;
  ram[12604]  = 1;
  ram[12605]  = 1;
  ram[12606]  = 1;
  ram[12607]  = 1;
  ram[12608]  = 1;
  ram[12609]  = 1;
  ram[12610]  = 1;
  ram[12611]  = 1;
  ram[12612]  = 1;
  ram[12613]  = 1;
  ram[12614]  = 1;
  ram[12615]  = 1;
  ram[12616]  = 1;
  ram[12617]  = 1;
  ram[12618]  = 1;
  ram[12619]  = 1;
  ram[12620]  = 1;
  ram[12621]  = 1;
  ram[12622]  = 1;
  ram[12623]  = 1;
  ram[12624]  = 1;
  ram[12625]  = 1;
  ram[12626]  = 1;
  ram[12627]  = 1;
  ram[12628]  = 1;
  ram[12629]  = 1;
  ram[12630]  = 0;
  ram[12631]  = 0;
  ram[12632]  = 0;
  ram[12633]  = 0;
  ram[12634]  = 0;
  ram[12635]  = 1;
  ram[12636]  = 1;
  ram[12637]  = 1;
  ram[12638]  = 1;
  ram[12639]  = 1;
  ram[12640]  = 1;
  ram[12641]  = 1;
  ram[12642]  = 1;
  ram[12643]  = 1;
  ram[12644]  = 1;
  ram[12645]  = 1;
  ram[12646]  = 1;
  ram[12647]  = 1;
  ram[12648]  = 0;
  ram[12649]  = 0;
  ram[12650]  = 0;
  ram[12651]  = 0;
  ram[12652]  = 1;
  ram[12653]  = 1;
  ram[12654]  = 1;
  ram[12655]  = 1;
  ram[12656]  = 1;
  ram[12657]  = 1;
  ram[12658]  = 1;
  ram[12659]  = 1;
  ram[12660]  = 1;
  ram[12661]  = 1;
  ram[12662]  = 1;
  ram[12663]  = 1;
  ram[12664]  = 1;
  ram[12665]  = 1;
  ram[12666]  = 1;
  ram[12667]  = 0;
  ram[12668]  = 0;
  ram[12669]  = 0;
  ram[12670]  = 0;
  ram[12671]  = 0;
  ram[12672]  = 1;
  ram[12673]  = 1;
  ram[12674]  = 1;
  ram[12675]  = 1;
  ram[12676]  = 1;
  ram[12677]  = 1;
  ram[12678]  = 1;
  ram[12679]  = 1;
  ram[12680]  = 1;
  ram[12681]  = 1;
  ram[12682]  = 1;
  ram[12683]  = 1;
  ram[12684]  = 1;
  ram[12685]  = 1;
  ram[12686]  = 1;
  ram[12687]  = 1;
  ram[12688]  = 1;
  ram[12689]  = 1;
  ram[12690]  = 1;
  ram[12691]  = 1;
  ram[12692]  = 1;
  ram[12693]  = 1;
  ram[12694]  = 1;
  ram[12695]  = 1;
  ram[12696]  = 1;
  ram[12697]  = 1;
  ram[12698]  = 1;
  ram[12699]  = 1;
  ram[12700]  = 1;
  ram[12701]  = 1;
  ram[12702]  = 1;
  ram[12703]  = 1;
  ram[12704]  = 1;
  ram[12705]  = 1;
  ram[12706]  = 1;
  ram[12707]  = 1;
  ram[12708]  = 1;
  ram[12709]  = 1;
  ram[12710]  = 1;
  ram[12711]  = 1;
  ram[12712]  = 1;
  ram[12713]  = 1;
  ram[12714]  = 1;
  ram[12715]  = 1;
  ram[12716]  = 1;
  ram[12717]  = 1;
  ram[12718]  = 1;
  ram[12719]  = 1;
  ram[12720]  = 1;
  ram[12721]  = 0;
  ram[12722]  = 0;
  ram[12723]  = 1;
  ram[12724]  = 1;
  ram[12725]  = 1;
  ram[12726]  = 1;
  ram[12727]  = 1;
  ram[12728]  = 0;
  ram[12729]  = 0;
  ram[12730]  = 1;
  ram[12731]  = 1;
  ram[12732]  = 0;
  ram[12733]  = 0;
  ram[12734]  = 0;
  ram[12735]  = 0;
  ram[12736]  = 1;
  ram[12737]  = 1;
  ram[12738]  = 1;
  ram[12739]  = 1;
  ram[12740]  = 1;
  ram[12741]  = 0;
  ram[12742]  = 0;
  ram[12743]  = 0;
  ram[12744]  = 0;
  ram[12745]  = 0;
  ram[12746]  = 0;
  ram[12747]  = 1;
  ram[12748]  = 1;
  ram[12749]  = 1;
  ram[12750]  = 1;
  ram[12751]  = 1;
  ram[12752]  = 1;
  ram[12753]  = 1;
  ram[12754]  = 1;
  ram[12755]  = 1;
  ram[12756]  = 1;
  ram[12757]  = 1;
  ram[12758]  = 1;
  ram[12759]  = 1;
  ram[12760]  = 1;
  ram[12761]  = 1;
  ram[12762]  = 1;
  ram[12763]  = 0;
  ram[12764]  = 0;
  ram[12765]  = 0;
  ram[12766]  = 1;
  ram[12767]  = 1;
  ram[12768]  = 1;
  ram[12769]  = 1;
  ram[12770]  = 1;
  ram[12771]  = 1;
  ram[12772]  = 1;
  ram[12773]  = 1;
  ram[12774]  = 1;
  ram[12775]  = 1;
  ram[12776]  = 1;
  ram[12777]  = 1;
  ram[12778]  = 1;
  ram[12779]  = 1;
  ram[12780]  = 1;
  ram[12781]  = 1;
  ram[12782]  = 1;
  ram[12783]  = 1;
  ram[12784]  = 1;
  ram[12785]  = 1;
  ram[12786]  = 1;
  ram[12787]  = 1;
  ram[12788]  = 1;
  ram[12789]  = 1;
  ram[12790]  = 1;
  ram[12791]  = 1;
  ram[12792]  = 1;
  ram[12793]  = 1;
  ram[12794]  = 1;
  ram[12795]  = 1;
  ram[12796]  = 1;
  ram[12797]  = 1;
  ram[12798]  = 1;
  ram[12799]  = 1;
  ram[12800]  = 1;
  ram[12801]  = 1;
  ram[12802]  = 1;
  ram[12803]  = 1;
  ram[12804]  = 1;
  ram[12805]  = 1;
  ram[12806]  = 1;
  ram[12807]  = 1;
  ram[12808]  = 1;
  ram[12809]  = 1;
  ram[12810]  = 1;
  ram[12811]  = 1;
  ram[12812]  = 1;
  ram[12813]  = 1;
  ram[12814]  = 1;
  ram[12815]  = 1;
  ram[12816]  = 1;
  ram[12817]  = 1;
  ram[12818]  = 1;
  ram[12819]  = 1;
  ram[12820]  = 1;
  ram[12821]  = 1;
  ram[12822]  = 1;
  ram[12823]  = 1;
  ram[12824]  = 1;
  ram[12825]  = 1;
  ram[12826]  = 1;
  ram[12827]  = 1;
  ram[12828]  = 1;
  ram[12829]  = 1;
  ram[12830]  = 1;
  ram[12831]  = 1;
  ram[12832]  = 1;
  ram[12833]  = 1;
  ram[12834]  = 1;
  ram[12835]  = 1;
  ram[12836]  = 1;
  ram[12837]  = 1;
  ram[12838]  = 1;
  ram[12839]  = 1;
  ram[12840]  = 1;
  ram[12841]  = 1;
  ram[12842]  = 1;
  ram[12843]  = 1;
  ram[12844]  = 1;
  ram[12845]  = 1;
  ram[12846]  = 1;
  ram[12847]  = 1;
  ram[12848]  = 1;
  ram[12849]  = 1;
  ram[12850]  = 1;
  ram[12851]  = 1;
  ram[12852]  = 1;
  ram[12853]  = 1;
  ram[12854]  = 1;
  ram[12855]  = 1;
  ram[12856]  = 1;
  ram[12857]  = 1;
  ram[12858]  = 1;
  ram[12859]  = 1;
  ram[12860]  = 1;
  ram[12861]  = 1;
  ram[12862]  = 1;
  ram[12863]  = 1;
  ram[12864]  = 1;
  ram[12865]  = 1;
  ram[12866]  = 1;
  ram[12867]  = 1;
  ram[12868]  = 1;
  ram[12869]  = 1;
  ram[12870]  = 1;
  ram[12871]  = 1;
  ram[12872]  = 1;
  ram[12873]  = 1;
  ram[12874]  = 1;
  ram[12875]  = 1;
  ram[12876]  = 1;
  ram[12877]  = 1;
  ram[12878]  = 1;
  ram[12879]  = 1;
  ram[12880]  = 1;
  ram[12881]  = 1;
  ram[12882]  = 1;
  ram[12883]  = 1;
  ram[12884]  = 1;
  ram[12885]  = 1;
  ram[12886]  = 1;
  ram[12887]  = 1;
  ram[12888]  = 1;
  ram[12889]  = 1;
  ram[12890]  = 1;
  ram[12891]  = 1;
  ram[12892]  = 1;
  ram[12893]  = 1;
  ram[12894]  = 1;
  ram[12895]  = 1;
  ram[12896]  = 1;
  ram[12897]  = 1;
  ram[12898]  = 1;
  ram[12899]  = 1;
  ram[12900]  = 1;
  ram[12901]  = 1;
  ram[12902]  = 1;
  ram[12903]  = 1;
  ram[12904]  = 1;
  ram[12905]  = 1;
  ram[12906]  = 1;
  ram[12907]  = 1;
  ram[12908]  = 1;
  ram[12909]  = 1;
  ram[12910]  = 1;
  ram[12911]  = 1;
  ram[12912]  = 1;
  ram[12913]  = 1;
  ram[12914]  = 1;
  ram[12915]  = 1;
  ram[12916]  = 1;
  ram[12917]  = 1;
  ram[12918]  = 1;
  ram[12919]  = 1;
  ram[12920]  = 1;
  ram[12921]  = 0;
  ram[12922]  = 0;
  ram[12923]  = 1;
  ram[12924]  = 1;
  ram[12925]  = 1;
  ram[12926]  = 1;
  ram[12927]  = 1;
  ram[12928]  = 0;
  ram[12929]  = 0;
  ram[12930]  = 1;
  ram[12931]  = 1;
  ram[12932]  = 1;
  ram[12933]  = 1;
  ram[12934]  = 1;
  ram[12935]  = 1;
  ram[12936]  = 1;
  ram[12937]  = 1;
  ram[12938]  = 1;
  ram[12939]  = 1;
  ram[12940]  = 1;
  ram[12941]  = 1;
  ram[12942]  = 1;
  ram[12943]  = 1;
  ram[12944]  = 1;
  ram[12945]  = 1;
  ram[12946]  = 1;
  ram[12947]  = 1;
  ram[12948]  = 1;
  ram[12949]  = 1;
  ram[12950]  = 1;
  ram[12951]  = 1;
  ram[12952]  = 1;
  ram[12953]  = 1;
  ram[12954]  = 1;
  ram[12955]  = 1;
  ram[12956]  = 1;
  ram[12957]  = 1;
  ram[12958]  = 1;
  ram[12959]  = 1;
  ram[12960]  = 1;
  ram[12961]  = 1;
  ram[12962]  = 1;
  ram[12963]  = 1;
  ram[12964]  = 1;
  ram[12965]  = 1;
  ram[12966]  = 1;
  ram[12967]  = 1;
  ram[12968]  = 1;
  ram[12969]  = 1;
  ram[12970]  = 1;
  ram[12971]  = 1;
  ram[12972]  = 1;
  ram[12973]  = 1;
  ram[12974]  = 1;
  ram[12975]  = 1;
  ram[12976]  = 1;
  ram[12977]  = 1;
  ram[12978]  = 1;
  ram[12979]  = 1;
  ram[12980]  = 1;
  ram[12981]  = 1;
  ram[12982]  = 1;
  ram[12983]  = 1;
  ram[12984]  = 1;
  ram[12985]  = 1;
  ram[12986]  = 1;
  ram[12987]  = 1;
  ram[12988]  = 1;
  ram[12989]  = 1;
  ram[12990]  = 1;
  ram[12991]  = 1;
  ram[12992]  = 1;
  ram[12993]  = 1;
  ram[12994]  = 1;
  ram[12995]  = 1;
  ram[12996]  = 1;
  ram[12997]  = 1;
  ram[12998]  = 1;
  ram[12999]  = 1;
  ram[13000]  = 1;
  ram[13001]  = 1;
  ram[13002]  = 1;
  ram[13003]  = 1;
  ram[13004]  = 1;
  ram[13005]  = 1;
  ram[13006]  = 1;
  ram[13007]  = 1;
  ram[13008]  = 1;
  ram[13009]  = 1;
  ram[13010]  = 1;
  ram[13011]  = 1;
  ram[13012]  = 1;
  ram[13013]  = 1;
  ram[13014]  = 1;
  ram[13015]  = 1;
  ram[13016]  = 1;
  ram[13017]  = 1;
  ram[13018]  = 1;
  ram[13019]  = 1;
  ram[13020]  = 1;
  ram[13021]  = 1;
  ram[13022]  = 1;
  ram[13023]  = 1;
  ram[13024]  = 1;
  ram[13025]  = 1;
  ram[13026]  = 1;
  ram[13027]  = 1;
  ram[13028]  = 1;
  ram[13029]  = 1;
  ram[13030]  = 1;
  ram[13031]  = 1;
  ram[13032]  = 1;
  ram[13033]  = 1;
  ram[13034]  = 1;
  ram[13035]  = 1;
  ram[13036]  = 1;
  ram[13037]  = 1;
  ram[13038]  = 1;
  ram[13039]  = 1;
  ram[13040]  = 1;
  ram[13041]  = 1;
  ram[13042]  = 1;
  ram[13043]  = 1;
  ram[13044]  = 1;
  ram[13045]  = 1;
  ram[13046]  = 1;
  ram[13047]  = 1;
  ram[13048]  = 1;
  ram[13049]  = 1;
  ram[13050]  = 1;
  ram[13051]  = 1;
  ram[13052]  = 1;
  ram[13053]  = 1;
  ram[13054]  = 1;
  ram[13055]  = 1;
  ram[13056]  = 1;
  ram[13057]  = 1;
  ram[13058]  = 1;
  ram[13059]  = 1;
  ram[13060]  = 1;
  ram[13061]  = 1;
  ram[13062]  = 1;
  ram[13063]  = 1;
  ram[13064]  = 1;
  ram[13065]  = 1;
  ram[13066]  = 1;
  ram[13067]  = 1;
  ram[13068]  = 1;
  ram[13069]  = 1;
  ram[13070]  = 1;
  ram[13071]  = 1;
  ram[13072]  = 1;
  ram[13073]  = 1;
  ram[13074]  = 1;
  ram[13075]  = 1;
  ram[13076]  = 1;
  ram[13077]  = 1;
  ram[13078]  = 1;
  ram[13079]  = 1;
  ram[13080]  = 1;
  ram[13081]  = 1;
  ram[13082]  = 1;
  ram[13083]  = 1;
  ram[13084]  = 1;
  ram[13085]  = 1;
  ram[13086]  = 1;
  ram[13087]  = 1;
  ram[13088]  = 1;
  ram[13089]  = 1;
  ram[13090]  = 1;
  ram[13091]  = 1;
  ram[13092]  = 1;
  ram[13093]  = 1;
  ram[13094]  = 1;
  ram[13095]  = 1;
  ram[13096]  = 1;
  ram[13097]  = 1;
  ram[13098]  = 1;
  ram[13099]  = 1;
  ram[13100]  = 1;
  ram[13101]  = 1;
  ram[13102]  = 1;
  ram[13103]  = 1;
  ram[13104]  = 1;
  ram[13105]  = 1;
  ram[13106]  = 1;
  ram[13107]  = 1;
  ram[13108]  = 1;
  ram[13109]  = 1;
  ram[13110]  = 1;
  ram[13111]  = 1;
  ram[13112]  = 1;
  ram[13113]  = 1;
  ram[13114]  = 1;
  ram[13115]  = 1;
  ram[13116]  = 1;
  ram[13117]  = 1;
  ram[13118]  = 1;
  ram[13119]  = 1;
  ram[13120]  = 1;
  ram[13121]  = 1;
  ram[13122]  = 1;
  ram[13123]  = 1;
  ram[13124]  = 1;
  ram[13125]  = 1;
  ram[13126]  = 1;
  ram[13127]  = 1;
  ram[13128]  = 1;
  ram[13129]  = 1;
  ram[13130]  = 1;
  ram[13131]  = 1;
  ram[13132]  = 1;
  ram[13133]  = 1;
  ram[13134]  = 1;
  ram[13135]  = 1;
  ram[13136]  = 1;
  ram[13137]  = 1;
  ram[13138]  = 1;
  ram[13139]  = 1;
  ram[13140]  = 1;
  ram[13141]  = 1;
  ram[13142]  = 1;
  ram[13143]  = 1;
  ram[13144]  = 1;
  ram[13145]  = 1;
  ram[13146]  = 1;
  ram[13147]  = 1;
  ram[13148]  = 1;
  ram[13149]  = 1;
  ram[13150]  = 1;
  ram[13151]  = 1;
  ram[13152]  = 1;
  ram[13153]  = 1;
  ram[13154]  = 1;
  ram[13155]  = 1;
  ram[13156]  = 1;
  ram[13157]  = 1;
  ram[13158]  = 1;
  ram[13159]  = 1;
  ram[13160]  = 1;
  ram[13161]  = 1;
  ram[13162]  = 1;
  ram[13163]  = 1;
  ram[13164]  = 1;
  ram[13165]  = 1;
  ram[13166]  = 1;
  ram[13167]  = 1;
  ram[13168]  = 1;
  ram[13169]  = 1;
  ram[13170]  = 1;
  ram[13171]  = 1;
  ram[13172]  = 1;
  ram[13173]  = 1;
  ram[13174]  = 1;
  ram[13175]  = 1;
  ram[13176]  = 1;
  ram[13177]  = 1;
  ram[13178]  = 1;
  ram[13179]  = 1;
  ram[13180]  = 1;
  ram[13181]  = 1;
  ram[13182]  = 1;
  ram[13183]  = 1;
  ram[13184]  = 1;
  ram[13185]  = 1;
  ram[13186]  = 1;
  ram[13187]  = 1;
  ram[13188]  = 1;
  ram[13189]  = 1;
  ram[13190]  = 1;
  ram[13191]  = 1;
  ram[13192]  = 1;
  ram[13193]  = 1;
  ram[13194]  = 1;
  ram[13195]  = 1;
  ram[13196]  = 1;
  ram[13197]  = 1;
  ram[13198]  = 1;
  ram[13199]  = 1;
  ram[13200]  = 1;
  ram[13201]  = 1;
  ram[13202]  = 1;
  ram[13203]  = 1;
  ram[13204]  = 1;
  ram[13205]  = 1;
  ram[13206]  = 1;
  ram[13207]  = 1;
  ram[13208]  = 1;
  ram[13209]  = 1;
  ram[13210]  = 1;
  ram[13211]  = 1;
  ram[13212]  = 1;
  ram[13213]  = 1;
  ram[13214]  = 1;
  ram[13215]  = 1;
  ram[13216]  = 1;
  ram[13217]  = 1;
  ram[13218]  = 1;
  ram[13219]  = 1;
  ram[13220]  = 1;
  ram[13221]  = 1;
  ram[13222]  = 1;
  ram[13223]  = 1;
  ram[13224]  = 1;
  ram[13225]  = 1;
  ram[13226]  = 1;
  ram[13227]  = 1;
  ram[13228]  = 1;
  ram[13229]  = 1;
  ram[13230]  = 1;
  ram[13231]  = 1;
  ram[13232]  = 1;
  ram[13233]  = 1;
  ram[13234]  = 1;
  ram[13235]  = 1;
  ram[13236]  = 1;
  ram[13237]  = 1;
  ram[13238]  = 1;
  ram[13239]  = 1;
  ram[13240]  = 1;
  ram[13241]  = 1;
  ram[13242]  = 1;
  ram[13243]  = 1;
  ram[13244]  = 1;
  ram[13245]  = 1;
  ram[13246]  = 1;
  ram[13247]  = 1;
  ram[13248]  = 1;
  ram[13249]  = 1;
  ram[13250]  = 1;
  ram[13251]  = 1;
  ram[13252]  = 1;
  ram[13253]  = 1;
  ram[13254]  = 1;
  ram[13255]  = 1;
  ram[13256]  = 1;
  ram[13257]  = 1;
  ram[13258]  = 1;
  ram[13259]  = 1;
  ram[13260]  = 1;
  ram[13261]  = 1;
  ram[13262]  = 1;
  ram[13263]  = 1;
  ram[13264]  = 1;
  ram[13265]  = 1;
  ram[13266]  = 1;
  ram[13267]  = 1;
  ram[13268]  = 1;
  ram[13269]  = 1;
  ram[13270]  = 1;
  ram[13271]  = 1;
  ram[13272]  = 1;
  ram[13273]  = 1;
  ram[13274]  = 1;
  ram[13275]  = 1;
  ram[13276]  = 1;
  ram[13277]  = 1;
  ram[13278]  = 1;
  ram[13279]  = 1;
  ram[13280]  = 1;
  ram[13281]  = 1;
  ram[13282]  = 1;
  ram[13283]  = 1;
  ram[13284]  = 1;
  ram[13285]  = 1;
  ram[13286]  = 1;
  ram[13287]  = 1;
  ram[13288]  = 1;
  ram[13289]  = 1;
  ram[13290]  = 1;
  ram[13291]  = 1;
  ram[13292]  = 1;
  ram[13293]  = 1;
  ram[13294]  = 1;
  ram[13295]  = 1;
  ram[13296]  = 1;
  ram[13297]  = 1;
  ram[13298]  = 1;
  ram[13299]  = 1;
  ram[13300]  = 1;
  ram[13301]  = 1;
  ram[13302]  = 1;
  ram[13303]  = 1;
  ram[13304]  = 1;
  ram[13305]  = 1;
  ram[13306]  = 1;
  ram[13307]  = 1;
  ram[13308]  = 1;
  ram[13309]  = 1;
  ram[13310]  = 1;
  ram[13311]  = 1;
  ram[13312]  = 1;
  ram[13313]  = 1;
  ram[13314]  = 1;
  ram[13315]  = 1;
  ram[13316]  = 1;
  ram[13317]  = 1;
  ram[13318]  = 1;
  ram[13319]  = 1;
  ram[13320]  = 1;
  ram[13321]  = 1;
  ram[13322]  = 1;
  ram[13323]  = 1;
  ram[13324]  = 1;
  ram[13325]  = 1;
  ram[13326]  = 1;
  ram[13327]  = 1;
  ram[13328]  = 1;
  ram[13329]  = 1;
  ram[13330]  = 1;
  ram[13331]  = 1;
  ram[13332]  = 1;
  ram[13333]  = 1;
  ram[13334]  = 1;
  ram[13335]  = 1;
  ram[13336]  = 1;
  ram[13337]  = 1;
  ram[13338]  = 1;
  ram[13339]  = 1;
  ram[13340]  = 1;
  ram[13341]  = 1;
  ram[13342]  = 1;
  ram[13343]  = 1;
  ram[13344]  = 1;
  ram[13345]  = 1;
  ram[13346]  = 1;
  ram[13347]  = 1;
  ram[13348]  = 1;
  ram[13349]  = 1;
  ram[13350]  = 1;
  ram[13351]  = 1;
  ram[13352]  = 1;
  ram[13353]  = 1;
  ram[13354]  = 1;
  ram[13355]  = 1;
  ram[13356]  = 1;
  ram[13357]  = 1;
  ram[13358]  = 1;
  ram[13359]  = 1;
  ram[13360]  = 1;
  ram[13361]  = 1;
  ram[13362]  = 1;
  ram[13363]  = 1;
  ram[13364]  = 1;
  ram[13365]  = 1;
  ram[13366]  = 1;
  ram[13367]  = 1;
  ram[13368]  = 1;
  ram[13369]  = 1;
  ram[13370]  = 1;
  ram[13371]  = 1;
  ram[13372]  = 1;
  ram[13373]  = 1;
  ram[13374]  = 1;
  ram[13375]  = 1;
  ram[13376]  = 1;
  ram[13377]  = 1;
  ram[13378]  = 1;
  ram[13379]  = 1;
  ram[13380]  = 1;
  ram[13381]  = 1;
  ram[13382]  = 1;
  ram[13383]  = 1;
  ram[13384]  = 1;
  ram[13385]  = 1;
  ram[13386]  = 1;
  ram[13387]  = 1;
  ram[13388]  = 1;
  ram[13389]  = 1;
  ram[13390]  = 1;
  ram[13391]  = 1;
  ram[13392]  = 1;
  ram[13393]  = 1;
  ram[13394]  = 1;
  ram[13395]  = 1;
  ram[13396]  = 1;
  ram[13397]  = 1;
  ram[13398]  = 1;
  ram[13399]  = 1;
  ram[13400]  = 1;
  ram[13401]  = 1;
  ram[13402]  = 1;
  ram[13403]  = 1;
  ram[13404]  = 1;
  ram[13405]  = 1;
  ram[13406]  = 1;
  ram[13407]  = 1;
  ram[13408]  = 1;
  ram[13409]  = 1;
  ram[13410]  = 1;
  ram[13411]  = 1;
  ram[13412]  = 1;
  ram[13413]  = 1;
  ram[13414]  = 1;
  ram[13415]  = 1;
  ram[13416]  = 1;
  ram[13417]  = 1;
  ram[13418]  = 1;
  ram[13419]  = 1;
  ram[13420]  = 1;
  ram[13421]  = 1;
  ram[13422]  = 1;
  ram[13423]  = 1;
  ram[13424]  = 1;
  ram[13425]  = 1;
  ram[13426]  = 1;
  ram[13427]  = 1;
  ram[13428]  = 1;
  ram[13429]  = 1;
  ram[13430]  = 1;
  ram[13431]  = 1;
  ram[13432]  = 1;
  ram[13433]  = 1;
  ram[13434]  = 1;
  ram[13435]  = 1;
  ram[13436]  = 1;
  ram[13437]  = 1;
  ram[13438]  = 1;
  ram[13439]  = 1;
  ram[13440]  = 1;
  ram[13441]  = 1;
  ram[13442]  = 1;
  ram[13443]  = 1;
  ram[13444]  = 1;
  ram[13445]  = 1;
  ram[13446]  = 1;
  ram[13447]  = 1;
  ram[13448]  = 1;
  ram[13449]  = 1;
  ram[13450]  = 1;
  ram[13451]  = 1;
  ram[13452]  = 1;
  ram[13453]  = 1;
  ram[13454]  = 1;
  ram[13455]  = 1;
  ram[13456]  = 1;
  ram[13457]  = 1;
  ram[13458]  = 1;
  ram[13459]  = 1;
  ram[13460]  = 1;
  ram[13461]  = 1;
  ram[13462]  = 1;
  ram[13463]  = 1;
  ram[13464]  = 1;
  ram[13465]  = 1;
  ram[13466]  = 1;
  ram[13467]  = 1;
  ram[13468]  = 1;
  ram[13469]  = 1;
  ram[13470]  = 1;
  ram[13471]  = 1;
  ram[13472]  = 1;
  ram[13473]  = 1;
  ram[13474]  = 1;
  ram[13475]  = 1;
  ram[13476]  = 1;
  ram[13477]  = 1;
  ram[13478]  = 1;
  ram[13479]  = 1;
  ram[13480]  = 1;
  ram[13481]  = 1;
  ram[13482]  = 1;
  ram[13483]  = 1;
  ram[13484]  = 1;
  ram[13485]  = 1;
  ram[13486]  = 1;
  ram[13487]  = 1;
  ram[13488]  = 1;
  ram[13489]  = 1;
  ram[13490]  = 1;
  ram[13491]  = 1;
  ram[13492]  = 1;
  ram[13493]  = 1;
  ram[13494]  = 1;
  ram[13495]  = 1;
  ram[13496]  = 1;
  ram[13497]  = 1;
  ram[13498]  = 1;
  ram[13499]  = 1;
  ram[13500]  = 1;
  ram[13501]  = 1;
  ram[13502]  = 1;
  ram[13503]  = 1;
  ram[13504]  = 1;
  ram[13505]  = 1;
  ram[13506]  = 1;
  ram[13507]  = 1;
  ram[13508]  = 1;
  ram[13509]  = 1;
  ram[13510]  = 1;
  ram[13511]  = 1;
  ram[13512]  = 1;
  ram[13513]  = 1;
  ram[13514]  = 1;
  ram[13515]  = 1;
  ram[13516]  = 1;
  ram[13517]  = 1;
  ram[13518]  = 1;
  ram[13519]  = 1;
  ram[13520]  = 1;
  ram[13521]  = 1;
  ram[13522]  = 1;
  ram[13523]  = 1;
  ram[13524]  = 1;
  ram[13525]  = 1;
  ram[13526]  = 1;
  ram[13527]  = 1;
  ram[13528]  = 1;
  ram[13529]  = 1;
  ram[13530]  = 1;
  ram[13531]  = 1;
  ram[13532]  = 1;
  ram[13533]  = 1;
  ram[13534]  = 1;
  ram[13535]  = 1;
  ram[13536]  = 1;
  ram[13537]  = 1;
  ram[13538]  = 1;
  ram[13539]  = 1;
  ram[13540]  = 1;
  ram[13541]  = 1;
  ram[13542]  = 1;
  ram[13543]  = 1;
  ram[13544]  = 1;
  ram[13545]  = 1;
  ram[13546]  = 1;
  ram[13547]  = 1;
  ram[13548]  = 1;
  ram[13549]  = 1;
  ram[13550]  = 1;
  ram[13551]  = 1;
  ram[13552]  = 1;
  ram[13553]  = 1;
  ram[13554]  = 1;
  ram[13555]  = 1;
  ram[13556]  = 1;
  ram[13557]  = 1;
  ram[13558]  = 1;
  ram[13559]  = 1;
  ram[13560]  = 1;
  ram[13561]  = 1;
  ram[13562]  = 1;
  ram[13563]  = 1;
  ram[13564]  = 1;
  ram[13565]  = 1;
  ram[13566]  = 1;
  ram[13567]  = 1;
  ram[13568]  = 1;
  ram[13569]  = 1;
  ram[13570]  = 1;
  ram[13571]  = 1;
  ram[13572]  = 1;
  ram[13573]  = 1;
  ram[13574]  = 1;
  ram[13575]  = 1;
  ram[13576]  = 1;
  ram[13577]  = 1;
  ram[13578]  = 1;
  ram[13579]  = 1;
  ram[13580]  = 1;
  ram[13581]  = 1;
  ram[13582]  = 1;
  ram[13583]  = 1;
  ram[13584]  = 1;
  ram[13585]  = 1;
  ram[13586]  = 1;
  ram[13587]  = 1;
  ram[13588]  = 1;
  ram[13589]  = 1;
  ram[13590]  = 1;
  ram[13591]  = 1;
  ram[13592]  = 1;
  ram[13593]  = 1;
  ram[13594]  = 1;
  ram[13595]  = 1;
  ram[13596]  = 1;
  ram[13597]  = 1;
  ram[13598]  = 1;
  ram[13599]  = 1;
  ram[13600]  = 1;
  ram[13601]  = 1;
  ram[13602]  = 1;
  ram[13603]  = 1;
  ram[13604]  = 1;
  ram[13605]  = 1;
  ram[13606]  = 1;
  ram[13607]  = 1;
  ram[13608]  = 1;
  ram[13609]  = 1;
  ram[13610]  = 1;
  ram[13611]  = 1;
  ram[13612]  = 1;
  ram[13613]  = 1;
  ram[13614]  = 1;
  ram[13615]  = 1;
  ram[13616]  = 1;
  ram[13617]  = 1;
  ram[13618]  = 1;
  ram[13619]  = 1;
  ram[13620]  = 1;
  ram[13621]  = 1;
  ram[13622]  = 1;
  ram[13623]  = 1;
  ram[13624]  = 1;
  ram[13625]  = 1;
  ram[13626]  = 1;
  ram[13627]  = 1;
  ram[13628]  = 1;
  ram[13629]  = 1;
  ram[13630]  = 1;
  ram[13631]  = 1;
  ram[13632]  = 1;
  ram[13633]  = 1;
  ram[13634]  = 1;
  ram[13635]  = 1;
  ram[13636]  = 1;
  ram[13637]  = 1;
  ram[13638]  = 1;
  ram[13639]  = 1;
  ram[13640]  = 1;
  ram[13641]  = 1;
  ram[13642]  = 1;
  ram[13643]  = 1;
  ram[13644]  = 1;
  ram[13645]  = 1;
  ram[13646]  = 1;
  ram[13647]  = 1;
  ram[13648]  = 1;
  ram[13649]  = 1;
  ram[13650]  = 1;
  ram[13651]  = 1;
  ram[13652]  = 1;
  ram[13653]  = 1;
  ram[13654]  = 1;
  ram[13655]  = 1;
  ram[13656]  = 1;
  ram[13657]  = 1;
  ram[13658]  = 1;
  ram[13659]  = 1;
  ram[13660]  = 1;
  ram[13661]  = 1;
  ram[13662]  = 1;
  ram[13663]  = 1;
  ram[13664]  = 1;
  ram[13665]  = 1;
  ram[13666]  = 1;
  ram[13667]  = 1;
  ram[13668]  = 1;
  ram[13669]  = 1;
  ram[13670]  = 1;
  ram[13671]  = 1;
  ram[13672]  = 1;
  ram[13673]  = 1;
  ram[13674]  = 1;
  ram[13675]  = 1;
  ram[13676]  = 1;
  ram[13677]  = 1;
  ram[13678]  = 1;
  ram[13679]  = 1;
  ram[13680]  = 1;
  ram[13681]  = 1;
  ram[13682]  = 1;
  ram[13683]  = 1;
  ram[13684]  = 1;
  ram[13685]  = 1;
  ram[13686]  = 1;
  ram[13687]  = 1;
  ram[13688]  = 1;
  ram[13689]  = 1;
  ram[13690]  = 1;
  ram[13691]  = 1;
  ram[13692]  = 1;
  ram[13693]  = 1;
  ram[13694]  = 1;
  ram[13695]  = 1;
  ram[13696]  = 1;
  ram[13697]  = 1;
  ram[13698]  = 1;
  ram[13699]  = 1;
  ram[13700]  = 1;
  ram[13701]  = 1;
  ram[13702]  = 1;
  ram[13703]  = 1;
  ram[13704]  = 1;
  ram[13705]  = 1;
  ram[13706]  = 1;
  ram[13707]  = 1;
  ram[13708]  = 1;
  ram[13709]  = 1;
  ram[13710]  = 1;
  ram[13711]  = 1;
  ram[13712]  = 1;
  ram[13713]  = 1;
  ram[13714]  = 1;
  ram[13715]  = 1;
  ram[13716]  = 1;
  ram[13717]  = 1;
  ram[13718]  = 1;
  ram[13719]  = 1;
  ram[13720]  = 1;
  ram[13721]  = 1;
  ram[13722]  = 1;
  ram[13723]  = 1;
  ram[13724]  = 1;
  ram[13725]  = 1;
  ram[13726]  = 1;
  ram[13727]  = 1;
  ram[13728]  = 1;
  ram[13729]  = 1;
  ram[13730]  = 1;
  ram[13731]  = 1;
  ram[13732]  = 1;
  ram[13733]  = 1;
  ram[13734]  = 1;
  ram[13735]  = 1;
  ram[13736]  = 1;
  ram[13737]  = 1;
  ram[13738]  = 1;
  ram[13739]  = 1;
  ram[13740]  = 1;
  ram[13741]  = 1;
  ram[13742]  = 1;
  ram[13743]  = 1;
  ram[13744]  = 1;
  ram[13745]  = 1;
  ram[13746]  = 1;
  ram[13747]  = 1;
  ram[13748]  = 1;
  ram[13749]  = 1;
  ram[13750]  = 1;
  ram[13751]  = 1;
  ram[13752]  = 1;
  ram[13753]  = 1;
  ram[13754]  = 1;
  ram[13755]  = 1;
  ram[13756]  = 1;
  ram[13757]  = 1;
  ram[13758]  = 1;
  ram[13759]  = 1;
  ram[13760]  = 1;
  ram[13761]  = 1;
  ram[13762]  = 1;
  ram[13763]  = 1;
  ram[13764]  = 1;
  ram[13765]  = 1;
  ram[13766]  = 1;
  ram[13767]  = 1;
  ram[13768]  = 1;
  ram[13769]  = 1;
  ram[13770]  = 1;
  ram[13771]  = 1;
  ram[13772]  = 1;
  ram[13773]  = 1;
  ram[13774]  = 1;
  ram[13775]  = 1;
  ram[13776]  = 1;
  ram[13777]  = 1;
  ram[13778]  = 1;
  ram[13779]  = 1;
  ram[13780]  = 1;
  ram[13781]  = 1;
  ram[13782]  = 1;
  ram[13783]  = 1;
  ram[13784]  = 1;
  ram[13785]  = 1;
  ram[13786]  = 1;
  ram[13787]  = 1;
  ram[13788]  = 1;
  ram[13789]  = 1;
  ram[13790]  = 1;
  ram[13791]  = 1;
  ram[13792]  = 1;
  ram[13793]  = 1;
  ram[13794]  = 1;
  ram[13795]  = 1;
  ram[13796]  = 1;
  ram[13797]  = 1;
  ram[13798]  = 1;
  ram[13799]  = 1;
  ram[13800]  = 1;
  ram[13801]  = 1;
  ram[13802]  = 1;
  ram[13803]  = 1;
  ram[13804]  = 1;
  ram[13805]  = 1;
  ram[13806]  = 1;
  ram[13807]  = 1;
  ram[13808]  = 1;
  ram[13809]  = 1;
  ram[13810]  = 1;
  ram[13811]  = 1;
  ram[13812]  = 1;
  ram[13813]  = 1;
  ram[13814]  = 1;
  ram[13815]  = 1;
  ram[13816]  = 1;
  ram[13817]  = 1;
  ram[13818]  = 1;
  ram[13819]  = 1;
  ram[13820]  = 1;
  ram[13821]  = 1;
  ram[13822]  = 1;
  ram[13823]  = 1;
  ram[13824]  = 1;
  ram[13825]  = 1;
  ram[13826]  = 1;
  ram[13827]  = 1;
  ram[13828]  = 1;
  ram[13829]  = 1;
  ram[13830]  = 1;
  ram[13831]  = 1;
  ram[13832]  = 1;
  ram[13833]  = 1;
  ram[13834]  = 1;
  ram[13835]  = 1;
  ram[13836]  = 1;
  ram[13837]  = 1;
  ram[13838]  = 1;
  ram[13839]  = 1;
  ram[13840]  = 1;
  ram[13841]  = 1;
  ram[13842]  = 1;
  ram[13843]  = 1;
  ram[13844]  = 1;
  ram[13845]  = 1;
  ram[13846]  = 1;
  ram[13847]  = 1;
  ram[13848]  = 1;
  ram[13849]  = 1;
  ram[13850]  = 1;
  ram[13851]  = 1;
  ram[13852]  = 1;
  ram[13853]  = 1;
  ram[13854]  = 1;
  ram[13855]  = 1;
  ram[13856]  = 1;
  ram[13857]  = 1;
  ram[13858]  = 1;
  ram[13859]  = 1;
  ram[13860]  = 1;
  ram[13861]  = 1;
  ram[13862]  = 1;
  ram[13863]  = 1;
  ram[13864]  = 1;
  ram[13865]  = 1;
  ram[13866]  = 1;
  ram[13867]  = 1;
  ram[13868]  = 1;
  ram[13869]  = 1;
  ram[13870]  = 1;
  ram[13871]  = 1;
  ram[13872]  = 1;
  ram[13873]  = 1;
  ram[13874]  = 1;
  ram[13875]  = 1;
  ram[13876]  = 1;
  ram[13877]  = 1;
  ram[13878]  = 1;
  ram[13879]  = 1;
  ram[13880]  = 1;
  ram[13881]  = 1;
  ram[13882]  = 1;
  ram[13883]  = 1;
  ram[13884]  = 1;
  ram[13885]  = 1;
  ram[13886]  = 1;
  ram[13887]  = 1;
  ram[13888]  = 1;
  ram[13889]  = 1;
  ram[13890]  = 1;
  ram[13891]  = 1;
  ram[13892]  = 1;
  ram[13893]  = 1;
  ram[13894]  = 1;
  ram[13895]  = 1;
  ram[13896]  = 1;
  ram[13897]  = 1;
  ram[13898]  = 1;
  ram[13899]  = 1;
  ram[13900]  = 1;
  ram[13901]  = 1;
  ram[13902]  = 1;
  ram[13903]  = 1;
  ram[13904]  = 1;
  ram[13905]  = 1;
  ram[13906]  = 1;
  ram[13907]  = 1;
  ram[13908]  = 1;
  ram[13909]  = 1;
  ram[13910]  = 1;
  ram[13911]  = 1;
  ram[13912]  = 1;
  ram[13913]  = 1;
  ram[13914]  = 1;
  ram[13915]  = 1;
  ram[13916]  = 1;
  ram[13917]  = 1;
  ram[13918]  = 1;
  ram[13919]  = 1;
  ram[13920]  = 1;
  ram[13921]  = 1;
  ram[13922]  = 1;
  ram[13923]  = 1;
  ram[13924]  = 1;
  ram[13925]  = 1;
  ram[13926]  = 1;
  ram[13927]  = 1;
  ram[13928]  = 1;
  ram[13929]  = 1;
  ram[13930]  = 1;
  ram[13931]  = 1;
  ram[13932]  = 1;
  ram[13933]  = 1;
  ram[13934]  = 1;
  ram[13935]  = 1;
  ram[13936]  = 1;
  ram[13937]  = 1;
  ram[13938]  = 1;
  ram[13939]  = 1;
  ram[13940]  = 1;
  ram[13941]  = 1;
  ram[13942]  = 1;
  ram[13943]  = 1;
  ram[13944]  = 1;
  ram[13945]  = 1;
  ram[13946]  = 1;
  ram[13947]  = 1;
  ram[13948]  = 1;
  ram[13949]  = 1;
  ram[13950]  = 1;
  ram[13951]  = 1;
  ram[13952]  = 1;
  ram[13953]  = 1;
  ram[13954]  = 1;
  ram[13955]  = 1;
  ram[13956]  = 1;
  ram[13957]  = 1;
  ram[13958]  = 1;
  ram[13959]  = 1;
  ram[13960]  = 1;
  ram[13961]  = 1;
  ram[13962]  = 1;
  ram[13963]  = 1;
  ram[13964]  = 1;
  ram[13965]  = 1;
  ram[13966]  = 1;
  ram[13967]  = 1;
  ram[13968]  = 1;
  ram[13969]  = 1;
  ram[13970]  = 1;
  ram[13971]  = 1;
  ram[13972]  = 1;
  ram[13973]  = 1;
  ram[13974]  = 1;
  ram[13975]  = 1;
  ram[13976]  = 1;
  ram[13977]  = 1;
  ram[13978]  = 1;
  ram[13979]  = 1;
  ram[13980]  = 1;
  ram[13981]  = 1;
  ram[13982]  = 1;
  ram[13983]  = 1;
  ram[13984]  = 1;
  ram[13985]  = 1;
  ram[13986]  = 1;
  ram[13987]  = 1;
  ram[13988]  = 1;
  ram[13989]  = 1;
  ram[13990]  = 1;
  ram[13991]  = 1;
  ram[13992]  = 1;
  ram[13993]  = 1;
  ram[13994]  = 1;
  ram[13995]  = 1;
  ram[13996]  = 1;
  ram[13997]  = 1;
  ram[13998]  = 1;
  ram[13999]  = 1;
  ram[14000]  = 1;
  ram[14001]  = 1;
  ram[14002]  = 1;
  ram[14003]  = 1;
  ram[14004]  = 1;
  ram[14005]  = 1;
  ram[14006]  = 1;
  ram[14007]  = 1;
  ram[14008]  = 1;
  ram[14009]  = 1;
  ram[14010]  = 1;
  ram[14011]  = 1;
  ram[14012]  = 1;
  ram[14013]  = 1;
  ram[14014]  = 1;
  ram[14015]  = 1;
  ram[14016]  = 1;
  ram[14017]  = 1;
  ram[14018]  = 1;
  ram[14019]  = 1;
  ram[14020]  = 1;
  ram[14021]  = 1;
  ram[14022]  = 1;
  ram[14023]  = 1;
  ram[14024]  = 1;
  ram[14025]  = 1;
  ram[14026]  = 1;
  ram[14027]  = 1;
  ram[14028]  = 1;
  ram[14029]  = 1;
  ram[14030]  = 1;
  ram[14031]  = 1;
  ram[14032]  = 1;
  ram[14033]  = 1;
  ram[14034]  = 1;
  ram[14035]  = 1;
  ram[14036]  = 1;
  ram[14037]  = 1;
  ram[14038]  = 1;
  ram[14039]  = 1;
  ram[14040]  = 1;
  ram[14041]  = 1;
  ram[14042]  = 1;
  ram[14043]  = 1;
  ram[14044]  = 1;
  ram[14045]  = 1;
  ram[14046]  = 1;
  ram[14047]  = 1;
  ram[14048]  = 1;
  ram[14049]  = 1;
  ram[14050]  = 1;
  ram[14051]  = 1;
  ram[14052]  = 1;
  ram[14053]  = 1;
  ram[14054]  = 1;
  ram[14055]  = 1;
  ram[14056]  = 1;
  ram[14057]  = 1;
  ram[14058]  = 1;
  ram[14059]  = 1;
  ram[14060]  = 1;
  ram[14061]  = 1;
  ram[14062]  = 1;
  ram[14063]  = 1;
  ram[14064]  = 1;
  ram[14065]  = 1;
  ram[14066]  = 1;
  ram[14067]  = 1;
  ram[14068]  = 1;
  ram[14069]  = 1;
  ram[14070]  = 1;
  ram[14071]  = 1;
  ram[14072]  = 1;
  ram[14073]  = 1;
  ram[14074]  = 1;
  ram[14075]  = 1;
  ram[14076]  = 1;
  ram[14077]  = 1;
  ram[14078]  = 1;
  ram[14079]  = 1;
  ram[14080]  = 1;
  ram[14081]  = 1;
  ram[14082]  = 1;
  ram[14083]  = 1;
  ram[14084]  = 1;
  ram[14085]  = 1;
  ram[14086]  = 1;
  ram[14087]  = 1;
  ram[14088]  = 1;
  ram[14089]  = 1;
  ram[14090]  = 1;
  ram[14091]  = 1;
  ram[14092]  = 1;
  ram[14093]  = 1;
  ram[14094]  = 1;
  ram[14095]  = 1;
  ram[14096]  = 1;
  ram[14097]  = 1;
  ram[14098]  = 1;
  ram[14099]  = 1;
  ram[14100]  = 1;
  ram[14101]  = 1;
  ram[14102]  = 1;
  ram[14103]  = 1;
  ram[14104]  = 1;
  ram[14105]  = 1;
  ram[14106]  = 1;
  ram[14107]  = 1;
  ram[14108]  = 1;
  ram[14109]  = 1;
  ram[14110]  = 1;
  ram[14111]  = 1;
  ram[14112]  = 1;
  ram[14113]  = 1;
  ram[14114]  = 1;
  ram[14115]  = 1;
  ram[14116]  = 1;
  ram[14117]  = 1;
  ram[14118]  = 1;
  ram[14119]  = 1;
  ram[14120]  = 1;
  ram[14121]  = 1;
  ram[14122]  = 1;
  ram[14123]  = 1;
  ram[14124]  = 1;
  ram[14125]  = 1;
  ram[14126]  = 1;
  ram[14127]  = 1;
  ram[14128]  = 1;
  ram[14129]  = 1;
  ram[14130]  = 1;
  ram[14131]  = 1;
  ram[14132]  = 1;
  ram[14133]  = 1;
  ram[14134]  = 1;
  ram[14135]  = 1;
  ram[14136]  = 1;
  ram[14137]  = 1;
  ram[14138]  = 1;
  ram[14139]  = 1;
  ram[14140]  = 1;
  ram[14141]  = 1;
  ram[14142]  = 1;
  ram[14143]  = 1;
  ram[14144]  = 1;
  ram[14145]  = 1;
  ram[14146]  = 1;
  ram[14147]  = 1;
  ram[14148]  = 1;
  ram[14149]  = 1;
  ram[14150]  = 1;
  ram[14151]  = 1;
  ram[14152]  = 1;
  ram[14153]  = 1;
  ram[14154]  = 1;
  ram[14155]  = 1;
  ram[14156]  = 1;
  ram[14157]  = 1;
  ram[14158]  = 1;
  ram[14159]  = 1;
  ram[14160]  = 1;
  ram[14161]  = 1;
  ram[14162]  = 1;
  ram[14163]  = 1;
  ram[14164]  = 1;
  ram[14165]  = 1;
  ram[14166]  = 1;
  ram[14167]  = 1;
  ram[14168]  = 1;
  ram[14169]  = 1;
  ram[14170]  = 1;
  ram[14171]  = 1;
  ram[14172]  = 1;
  ram[14173]  = 1;
  ram[14174]  = 1;
  ram[14175]  = 1;
  ram[14176]  = 1;
  ram[14177]  = 1;
  ram[14178]  = 1;
  ram[14179]  = 1;
  ram[14180]  = 1;
  ram[14181]  = 1;
  ram[14182]  = 1;
  ram[14183]  = 1;
  ram[14184]  = 1;
  ram[14185]  = 1;
  ram[14186]  = 1;
  ram[14187]  = 1;
  ram[14188]  = 1;
  ram[14189]  = 1;
  ram[14190]  = 1;
  ram[14191]  = 1;
  ram[14192]  = 1;
  ram[14193]  = 1;
  ram[14194]  = 1;
  ram[14195]  = 1;
  ram[14196]  = 1;
  ram[14197]  = 1;
  ram[14198]  = 1;
  ram[14199]  = 1;
  ram[14200]  = 1;
  ram[14201]  = 1;
  ram[14202]  = 1;
  ram[14203]  = 1;
  ram[14204]  = 1;
  ram[14205]  = 1;
  ram[14206]  = 1;
  ram[14207]  = 1;
  ram[14208]  = 1;
  ram[14209]  = 1;
  ram[14210]  = 1;
  ram[14211]  = 1;
  ram[14212]  = 1;
  ram[14213]  = 1;
  ram[14214]  = 1;
  ram[14215]  = 1;
  ram[14216]  = 1;
  ram[14217]  = 1;
  ram[14218]  = 1;
  ram[14219]  = 1;
  ram[14220]  = 1;
  ram[14221]  = 1;
  ram[14222]  = 1;
  ram[14223]  = 1;
  ram[14224]  = 1;
  ram[14225]  = 1;
  ram[14226]  = 1;
  ram[14227]  = 1;
  ram[14228]  = 1;
  ram[14229]  = 1;
  ram[14230]  = 1;
  ram[14231]  = 1;
  ram[14232]  = 1;
  ram[14233]  = 1;
  ram[14234]  = 1;
  ram[14235]  = 1;
  ram[14236]  = 1;
  ram[14237]  = 1;
  ram[14238]  = 1;
  ram[14239]  = 1;
  ram[14240]  = 1;
  ram[14241]  = 1;
  ram[14242]  = 1;
  ram[14243]  = 1;
  ram[14244]  = 1;
  ram[14245]  = 1;
  ram[14246]  = 1;
  ram[14247]  = 1;
  ram[14248]  = 1;
  ram[14249]  = 1;
  ram[14250]  = 1;
  ram[14251]  = 1;
  ram[14252]  = 1;
  ram[14253]  = 1;
  ram[14254]  = 1;
  ram[14255]  = 1;
  ram[14256]  = 1;
  ram[14257]  = 1;
  ram[14258]  = 1;
  ram[14259]  = 1;
  ram[14260]  = 1;
  ram[14261]  = 1;
  ram[14262]  = 1;
  ram[14263]  = 1;
  ram[14264]  = 1;
  ram[14265]  = 1;
  ram[14266]  = 1;
  ram[14267]  = 1;
  ram[14268]  = 1;
  ram[14269]  = 1;
  ram[14270]  = 1;
  ram[14271]  = 1;
  ram[14272]  = 1;
  ram[14273]  = 1;
  ram[14274]  = 1;
  ram[14275]  = 1;
  ram[14276]  = 1;
  ram[14277]  = 1;
  ram[14278]  = 1;
  ram[14279]  = 1;
  ram[14280]  = 1;
  ram[14281]  = 1;
  ram[14282]  = 1;
  ram[14283]  = 1;
  ram[14284]  = 1;
  ram[14285]  = 1;
  ram[14286]  = 1;
  ram[14287]  = 1;
  ram[14288]  = 1;
  ram[14289]  = 1;
  ram[14290]  = 1;
  ram[14291]  = 1;
  ram[14292]  = 1;
  ram[14293]  = 1;
  ram[14294]  = 1;
  ram[14295]  = 1;
  ram[14296]  = 1;
  ram[14297]  = 1;
  ram[14298]  = 1;
  ram[14299]  = 1;
  ram[14300]  = 1;
  ram[14301]  = 1;
  ram[14302]  = 1;
  ram[14303]  = 1;
  ram[14304]  = 1;
  ram[14305]  = 1;
  ram[14306]  = 1;
  ram[14307]  = 1;
  ram[14308]  = 1;
  ram[14309]  = 1;
  ram[14310]  = 1;
  ram[14311]  = 1;
  ram[14312]  = 1;
  ram[14313]  = 1;
  ram[14314]  = 1;
  ram[14315]  = 1;
  ram[14316]  = 1;
  ram[14317]  = 1;
  ram[14318]  = 1;
  ram[14319]  = 1;
  ram[14320]  = 1;
  ram[14321]  = 1;
  ram[14322]  = 1;
  ram[14323]  = 1;
  ram[14324]  = 1;
  ram[14325]  = 1;
  ram[14326]  = 1;
  ram[14327]  = 1;
  ram[14328]  = 1;
  ram[14329]  = 1;
  ram[14330]  = 1;
  ram[14331]  = 1;
  ram[14332]  = 1;
  ram[14333]  = 1;
  ram[14334]  = 1;
  ram[14335]  = 1;
  ram[14336]  = 1;
  ram[14337]  = 1;
  ram[14338]  = 1;
  ram[14339]  = 1;
  ram[14340]  = 1;
  ram[14341]  = 1;
  ram[14342]  = 1;
  ram[14343]  = 1;
  ram[14344]  = 1;
  ram[14345]  = 1;
  ram[14346]  = 1;
  ram[14347]  = 1;
  ram[14348]  = 1;
  ram[14349]  = 1;
  ram[14350]  = 1;
  ram[14351]  = 1;
  ram[14352]  = 1;
  ram[14353]  = 1;
  ram[14354]  = 1;
  ram[14355]  = 1;
  ram[14356]  = 1;
  ram[14357]  = 1;
  ram[14358]  = 1;
  ram[14359]  = 1;
  ram[14360]  = 1;
  ram[14361]  = 1;
  ram[14362]  = 1;
  ram[14363]  = 1;
  ram[14364]  = 1;
  ram[14365]  = 1;
  ram[14366]  = 1;
  ram[14367]  = 1;
  ram[14368]  = 1;
  ram[14369]  = 1;
  ram[14370]  = 1;
  ram[14371]  = 1;
  ram[14372]  = 1;
  ram[14373]  = 1;
  ram[14374]  = 1;
  ram[14375]  = 1;
  ram[14376]  = 1;
  ram[14377]  = 1;
  ram[14378]  = 1;
  ram[14379]  = 1;
  ram[14380]  = 1;
  ram[14381]  = 1;
  ram[14382]  = 1;
  ram[14383]  = 1;
  ram[14384]  = 1;
  ram[14385]  = 1;
  ram[14386]  = 1;
  ram[14387]  = 1;
  ram[14388]  = 1;
  ram[14389]  = 1;
  ram[14390]  = 1;
  ram[14391]  = 1;
  ram[14392]  = 1;
  ram[14393]  = 1;
  ram[14394]  = 1;
  ram[14395]  = 1;
  ram[14396]  = 1;
  ram[14397]  = 1;
  ram[14398]  = 1;
  ram[14399]  = 1;
  ram[14400]  = 1;
  ram[14401]  = 1;
  ram[14402]  = 1;
  ram[14403]  = 1;
  ram[14404]  = 1;
  ram[14405]  = 1;
  ram[14406]  = 1;
  ram[14407]  = 1;
  ram[14408]  = 1;
  ram[14409]  = 1;
  ram[14410]  = 1;
  ram[14411]  = 1;
  ram[14412]  = 1;
  ram[14413]  = 1;
  ram[14414]  = 1;
  ram[14415]  = 1;
  ram[14416]  = 1;
  ram[14417]  = 1;
  ram[14418]  = 1;
  ram[14419]  = 1;
  ram[14420]  = 1;
  ram[14421]  = 1;
  ram[14422]  = 1;
  ram[14423]  = 1;
  ram[14424]  = 1;
  ram[14425]  = 1;
  ram[14426]  = 1;
  ram[14427]  = 1;
  ram[14428]  = 1;
  ram[14429]  = 1;
  ram[14430]  = 1;
  ram[14431]  = 1;
  ram[14432]  = 1;
  ram[14433]  = 1;
  ram[14434]  = 1;
  ram[14435]  = 1;
  ram[14436]  = 1;
  ram[14437]  = 1;
  ram[14438]  = 1;
  ram[14439]  = 1;
  ram[14440]  = 1;
  ram[14441]  = 1;
  ram[14442]  = 1;
  ram[14443]  = 1;
  ram[14444]  = 1;
  ram[14445]  = 1;
  ram[14446]  = 1;
  ram[14447]  = 1;
  ram[14448]  = 1;
  ram[14449]  = 1;
  ram[14450]  = 1;
  ram[14451]  = 1;
  ram[14452]  = 1;
  ram[14453]  = 1;
  ram[14454]  = 1;
  ram[14455]  = 1;
  ram[14456]  = 1;
  ram[14457]  = 1;
  ram[14458]  = 1;
  ram[14459]  = 1;
  ram[14460]  = 1;
  ram[14461]  = 1;
  ram[14462]  = 1;
  ram[14463]  = 1;
  ram[14464]  = 1;
  ram[14465]  = 1;
  ram[14466]  = 1;
  ram[14467]  = 1;
  ram[14468]  = 1;
  ram[14469]  = 1;
  ram[14470]  = 1;
  ram[14471]  = 1;
  ram[14472]  = 1;
  ram[14473]  = 1;
  ram[14474]  = 1;
  ram[14475]  = 1;
  ram[14476]  = 1;
  ram[14477]  = 1;
  ram[14478]  = 1;
  ram[14479]  = 1;
  ram[14480]  = 1;
  ram[14481]  = 1;
  ram[14482]  = 1;
  ram[14483]  = 1;
  ram[14484]  = 1;
  ram[14485]  = 1;
  ram[14486]  = 1;
  ram[14487]  = 1;
  ram[14488]  = 1;
  ram[14489]  = 1;
  ram[14490]  = 1;
  ram[14491]  = 1;
  ram[14492]  = 1;
  ram[14493]  = 1;
  ram[14494]  = 1;
  ram[14495]  = 1;
  ram[14496]  = 1;
  ram[14497]  = 1;
  ram[14498]  = 1;
  ram[14499]  = 1;
  ram[14500]  = 1;
  ram[14501]  = 1;
  ram[14502]  = 1;
  ram[14503]  = 1;
  ram[14504]  = 1;
  ram[14505]  = 1;
  ram[14506]  = 1;
  ram[14507]  = 1;
  ram[14508]  = 1;
  ram[14509]  = 1;
  ram[14510]  = 1;
  ram[14511]  = 1;
  ram[14512]  = 1;
  ram[14513]  = 1;
  ram[14514]  = 1;
  ram[14515]  = 1;
  ram[14516]  = 1;
  ram[14517]  = 1;
  ram[14518]  = 1;
  ram[14519]  = 1;
  ram[14520]  = 1;
  ram[14521]  = 1;
  ram[14522]  = 1;
  ram[14523]  = 1;
  ram[14524]  = 1;
  ram[14525]  = 1;
  ram[14526]  = 1;
  ram[14527]  = 1;
  ram[14528]  = 1;
  ram[14529]  = 1;
  ram[14530]  = 1;
  ram[14531]  = 1;
  ram[14532]  = 1;
  ram[14533]  = 1;
  ram[14534]  = 1;
  ram[14535]  = 1;
  ram[14536]  = 1;
  ram[14537]  = 1;
  ram[14538]  = 1;
  ram[14539]  = 1;
  ram[14540]  = 1;
  ram[14541]  = 1;
  ram[14542]  = 1;
  ram[14543]  = 1;
  ram[14544]  = 1;
  ram[14545]  = 1;
  ram[14546]  = 1;
  ram[14547]  = 1;
  ram[14548]  = 1;
  ram[14549]  = 1;
  ram[14550]  = 1;
  ram[14551]  = 1;
  ram[14552]  = 1;
  ram[14553]  = 1;
  ram[14554]  = 1;
  ram[14555]  = 1;
  ram[14556]  = 1;
  ram[14557]  = 1;
  ram[14558]  = 1;
  ram[14559]  = 1;
  ram[14560]  = 1;
  ram[14561]  = 1;
  ram[14562]  = 1;
  ram[14563]  = 1;
  ram[14564]  = 1;
  ram[14565]  = 1;
  ram[14566]  = 1;
  ram[14567]  = 1;
  ram[14568]  = 1;
  ram[14569]  = 1;
  ram[14570]  = 1;
  ram[14571]  = 1;
  ram[14572]  = 1;
  ram[14573]  = 1;
  ram[14574]  = 1;
  ram[14575]  = 1;
  ram[14576]  = 1;
  ram[14577]  = 1;
  ram[14578]  = 1;
  ram[14579]  = 1;
  ram[14580]  = 1;
  ram[14581]  = 1;
  ram[14582]  = 1;
  ram[14583]  = 1;
  ram[14584]  = 1;
  ram[14585]  = 1;
  ram[14586]  = 1;
  ram[14587]  = 1;
  ram[14588]  = 1;
  ram[14589]  = 1;
  ram[14590]  = 1;
  ram[14591]  = 1;
  ram[14592]  = 1;
  ram[14593]  = 1;
  ram[14594]  = 1;
  ram[14595]  = 1;
  ram[14596]  = 1;
  ram[14597]  = 1;
  ram[14598]  = 1;
  ram[14599]  = 1;
  ram[14600]  = 1;
  ram[14601]  = 1;
  ram[14602]  = 1;
  ram[14603]  = 1;
  ram[14604]  = 1;
  ram[14605]  = 1;
  ram[14606]  = 1;
  ram[14607]  = 1;
  ram[14608]  = 1;
  ram[14609]  = 1;
  ram[14610]  = 1;
  ram[14611]  = 1;
  ram[14612]  = 1;
  ram[14613]  = 1;
  ram[14614]  = 1;
  ram[14615]  = 1;
  ram[14616]  = 1;
  ram[14617]  = 1;
  ram[14618]  = 1;
  ram[14619]  = 1;
  ram[14620]  = 1;
  ram[14621]  = 1;
  ram[14622]  = 1;
  ram[14623]  = 1;
  ram[14624]  = 1;
  ram[14625]  = 1;
  ram[14626]  = 1;
  ram[14627]  = 1;
  ram[14628]  = 1;
  ram[14629]  = 1;
  ram[14630]  = 1;
  ram[14631]  = 1;
  ram[14632]  = 1;
  ram[14633]  = 1;
  ram[14634]  = 1;
  ram[14635]  = 1;
  ram[14636]  = 1;
  ram[14637]  = 1;
  ram[14638]  = 1;
  ram[14639]  = 1;
  ram[14640]  = 1;
  ram[14641]  = 1;
  ram[14642]  = 1;
  ram[14643]  = 1;
  ram[14644]  = 1;
  ram[14645]  = 1;
  ram[14646]  = 1;
  ram[14647]  = 1;
  ram[14648]  = 1;
  ram[14649]  = 1;
  ram[14650]  = 1;
  ram[14651]  = 1;
  ram[14652]  = 1;
  ram[14653]  = 1;
  ram[14654]  = 1;
  ram[14655]  = 1;
  ram[14656]  = 1;
  ram[14657]  = 1;
  ram[14658]  = 1;
  ram[14659]  = 1;
  ram[14660]  = 1;
  ram[14661]  = 1;
  ram[14662]  = 1;
  ram[14663]  = 1;
  ram[14664]  = 1;
  ram[14665]  = 1;
  ram[14666]  = 1;
  ram[14667]  = 1;
  ram[14668]  = 1;
  ram[14669]  = 1;
  ram[14670]  = 1;
  ram[14671]  = 1;
  ram[14672]  = 1;
  ram[14673]  = 1;
  ram[14674]  = 1;
  ram[14675]  = 1;
  ram[14676]  = 1;
  ram[14677]  = 1;
  ram[14678]  = 1;
  ram[14679]  = 1;
  ram[14680]  = 1;
  ram[14681]  = 1;
  ram[14682]  = 1;
  ram[14683]  = 1;
  ram[14684]  = 1;
  ram[14685]  = 1;
  ram[14686]  = 1;
  ram[14687]  = 1;
  ram[14688]  = 1;
  ram[14689]  = 1;
  ram[14690]  = 1;
  ram[14691]  = 1;
  ram[14692]  = 1;
  ram[14693]  = 1;
  ram[14694]  = 1;
  ram[14695]  = 1;
  ram[14696]  = 1;
  ram[14697]  = 1;
  ram[14698]  = 1;
  ram[14699]  = 1;
  ram[14700]  = 1;
  ram[14701]  = 1;
  ram[14702]  = 1;
  ram[14703]  = 1;
  ram[14704]  = 1;
  ram[14705]  = 1;
  ram[14706]  = 1;
  ram[14707]  = 1;
  ram[14708]  = 1;
  ram[14709]  = 1;
  ram[14710]  = 1;
  ram[14711]  = 1;
  ram[14712]  = 1;
  ram[14713]  = 1;
  ram[14714]  = 1;
  ram[14715]  = 1;
  ram[14716]  = 1;
  ram[14717]  = 1;
  ram[14718]  = 1;
  ram[14719]  = 1;
  ram[14720]  = 1;
  ram[14721]  = 1;
  ram[14722]  = 1;
  ram[14723]  = 1;
  ram[14724]  = 1;
  ram[14725]  = 1;
  ram[14726]  = 1;
  ram[14727]  = 1;
  ram[14728]  = 1;
  ram[14729]  = 1;
  ram[14730]  = 1;
  ram[14731]  = 1;
  ram[14732]  = 1;
  ram[14733]  = 1;
  ram[14734]  = 1;
  ram[14735]  = 1;
  ram[14736]  = 1;
  ram[14737]  = 1;
  ram[14738]  = 1;
  ram[14739]  = 1;
  ram[14740]  = 1;
  ram[14741]  = 1;
  ram[14742]  = 1;
  ram[14743]  = 1;
  ram[14744]  = 1;
  ram[14745]  = 1;
  ram[14746]  = 1;
  ram[14747]  = 1;
  ram[14748]  = 1;
  ram[14749]  = 1;
  ram[14750]  = 1;
  ram[14751]  = 1;
  ram[14752]  = 1;
  ram[14753]  = 1;
  ram[14754]  = 1;
  ram[14755]  = 1;
  ram[14756]  = 1;
  ram[14757]  = 1;
  ram[14758]  = 1;
  ram[14759]  = 1;
  ram[14760]  = 1;
  ram[14761]  = 1;
  ram[14762]  = 1;
  ram[14763]  = 1;
  ram[14764]  = 1;
  ram[14765]  = 1;
  ram[14766]  = 1;
  ram[14767]  = 1;
  ram[14768]  = 1;
  ram[14769]  = 1;
  ram[14770]  = 1;
  ram[14771]  = 1;
  ram[14772]  = 1;
  ram[14773]  = 1;
  ram[14774]  = 1;
  ram[14775]  = 1;
  ram[14776]  = 1;
  ram[14777]  = 1;
  ram[14778]  = 1;
  ram[14779]  = 1;
  ram[14780]  = 1;
  ram[14781]  = 1;
  ram[14782]  = 1;
  ram[14783]  = 1;
  ram[14784]  = 1;
  ram[14785]  = 1;
  ram[14786]  = 1;
  ram[14787]  = 1;
  ram[14788]  = 1;
  ram[14789]  = 1;
  ram[14790]  = 1;
  ram[14791]  = 1;
  ram[14792]  = 1;
  ram[14793]  = 1;
  ram[14794]  = 1;
  ram[14795]  = 1;
  ram[14796]  = 1;
  ram[14797]  = 1;
  ram[14798]  = 1;
  ram[14799]  = 1;
  ram[14800]  = 1;
  ram[14801]  = 1;
  ram[14802]  = 1;
  ram[14803]  = 1;
  ram[14804]  = 1;
  ram[14805]  = 1;
  ram[14806]  = 1;
  ram[14807]  = 1;
  ram[14808]  = 1;
  ram[14809]  = 1;
  ram[14810]  = 1;
  ram[14811]  = 1;
  ram[14812]  = 1;
  ram[14813]  = 1;
  ram[14814]  = 1;
  ram[14815]  = 1;
  ram[14816]  = 1;
  ram[14817]  = 1;
  ram[14818]  = 1;
  ram[14819]  = 1;
  ram[14820]  = 1;
  ram[14821]  = 1;
  ram[14822]  = 1;
  ram[14823]  = 1;
  ram[14824]  = 1;
  ram[14825]  = 1;
  ram[14826]  = 1;
  ram[14827]  = 1;
  ram[14828]  = 1;
  ram[14829]  = 1;
  ram[14830]  = 1;
  ram[14831]  = 1;
  ram[14832]  = 1;
  ram[14833]  = 1;
  ram[14834]  = 1;
  ram[14835]  = 1;
  ram[14836]  = 1;
  ram[14837]  = 1;
  ram[14838]  = 1;
  ram[14839]  = 1;
  ram[14840]  = 1;
  ram[14841]  = 1;
  ram[14842]  = 1;
  ram[14843]  = 1;
  ram[14844]  = 1;
  ram[14845]  = 1;
  ram[14846]  = 1;
  ram[14847]  = 1;
  ram[14848]  = 1;
  ram[14849]  = 1;
  ram[14850]  = 1;
  ram[14851]  = 1;
  ram[14852]  = 1;
  ram[14853]  = 1;
  ram[14854]  = 1;
  ram[14855]  = 1;
  ram[14856]  = 1;
  ram[14857]  = 1;
  ram[14858]  = 1;
  ram[14859]  = 1;
  ram[14860]  = 1;
  ram[14861]  = 1;
  ram[14862]  = 1;
  ram[14863]  = 1;
  ram[14864]  = 1;
  ram[14865]  = 1;
  ram[14866]  = 1;
  ram[14867]  = 1;
  ram[14868]  = 1;
  ram[14869]  = 1;
  ram[14870]  = 1;
  ram[14871]  = 1;
  ram[14872]  = 1;
  ram[14873]  = 1;
  ram[14874]  = 1;
  ram[14875]  = 1;
  ram[14876]  = 1;
  ram[14877]  = 1;
  ram[14878]  = 1;
  ram[14879]  = 1;
  ram[14880]  = 1;
  ram[14881]  = 1;
  ram[14882]  = 1;
  ram[14883]  = 1;
  ram[14884]  = 1;
  ram[14885]  = 1;
  ram[14886]  = 1;
  ram[14887]  = 1;
  ram[14888]  = 1;
  ram[14889]  = 1;
  ram[14890]  = 1;
  ram[14891]  = 1;
  ram[14892]  = 1;
  ram[14893]  = 1;
  ram[14894]  = 1;
  ram[14895]  = 1;
  ram[14896]  = 1;
  ram[14897]  = 1;
  ram[14898]  = 1;
  ram[14899]  = 1;
  ram[14900]  = 1;
  ram[14901]  = 1;
  ram[14902]  = 1;
  ram[14903]  = 1;
  ram[14904]  = 1;
  ram[14905]  = 1;
  ram[14906]  = 1;
  ram[14907]  = 1;
  ram[14908]  = 1;
  ram[14909]  = 1;
  ram[14910]  = 1;
  ram[14911]  = 1;
  ram[14912]  = 1;
  ram[14913]  = 1;
  ram[14914]  = 1;
  ram[14915]  = 1;
  ram[14916]  = 1;
  ram[14917]  = 1;
  ram[14918]  = 1;
  ram[14919]  = 1;
  ram[14920]  = 1;
  ram[14921]  = 1;
  ram[14922]  = 1;
  ram[14923]  = 1;
  ram[14924]  = 1;
  ram[14925]  = 1;
  ram[14926]  = 1;
  ram[14927]  = 1;
  ram[14928]  = 1;
  ram[14929]  = 1;
  ram[14930]  = 1;
  ram[14931]  = 1;
  ram[14932]  = 1;
  ram[14933]  = 1;
  ram[14934]  = 1;
  ram[14935]  = 1;
  ram[14936]  = 1;
  ram[14937]  = 1;
  ram[14938]  = 1;
  ram[14939]  = 1;
  ram[14940]  = 1;
  ram[14941]  = 1;
  ram[14942]  = 1;
  ram[14943]  = 1;
  ram[14944]  = 1;
  ram[14945]  = 1;
  ram[14946]  = 1;
  ram[14947]  = 1;
  ram[14948]  = 1;
  ram[14949]  = 1;
  ram[14950]  = 1;
  ram[14951]  = 1;
  ram[14952]  = 1;
  ram[14953]  = 1;
  ram[14954]  = 1;
  ram[14955]  = 1;
  ram[14956]  = 1;
  ram[14957]  = 1;
  ram[14958]  = 1;
  ram[14959]  = 1;
  ram[14960]  = 1;
  ram[14961]  = 1;
  ram[14962]  = 1;
  ram[14963]  = 1;
  ram[14964]  = 1;
  ram[14965]  = 1;
  ram[14966]  = 1;
  ram[14967]  = 1;
  ram[14968]  = 1;
  ram[14969]  = 1;
  ram[14970]  = 1;
  ram[14971]  = 1;
  ram[14972]  = 1;
  ram[14973]  = 1;
  ram[14974]  = 1;
  ram[14975]  = 1;
  ram[14976]  = 1;
  ram[14977]  = 1;
  ram[14978]  = 1;
  ram[14979]  = 1;
  ram[14980]  = 1;
  ram[14981]  = 1;
  ram[14982]  = 1;
  ram[14983]  = 1;
  ram[14984]  = 1;
  ram[14985]  = 1;
  ram[14986]  = 1;
  ram[14987]  = 1;
  ram[14988]  = 1;
  ram[14989]  = 1;
  ram[14990]  = 1;
  ram[14991]  = 1;
  ram[14992]  = 1;
  ram[14993]  = 1;
  ram[14994]  = 1;
  ram[14995]  = 1;
  ram[14996]  = 1;
  ram[14997]  = 1;
  ram[14998]  = 1;
  ram[14999]  = 1;
  ram[15000]  = 1;
  ram[15001]  = 1;
  ram[15002]  = 1;
  ram[15003]  = 1;
  ram[15004]  = 1;
  ram[15005]  = 1;
  ram[15006]  = 1;
  ram[15007]  = 1;
  ram[15008]  = 1;
  ram[15009]  = 1;
  ram[15010]  = 1;
  ram[15011]  = 1;
  ram[15012]  = 1;
  ram[15013]  = 1;
  ram[15014]  = 1;
  ram[15015]  = 1;
  ram[15016]  = 1;
  ram[15017]  = 1;
  ram[15018]  = 1;
  ram[15019]  = 1;
  ram[15020]  = 1;
  ram[15021]  = 1;
  ram[15022]  = 1;
  ram[15023]  = 1;
  ram[15024]  = 1;
  ram[15025]  = 1;
  ram[15026]  = 1;
  ram[15027]  = 1;
  ram[15028]  = 1;
  ram[15029]  = 1;
  ram[15030]  = 1;
  ram[15031]  = 1;
  ram[15032]  = 1;
  ram[15033]  = 1;
  ram[15034]  = 1;
  ram[15035]  = 1;
  ram[15036]  = 1;
  ram[15037]  = 1;
  ram[15038]  = 1;
  ram[15039]  = 1;
  ram[15040]  = 1;
  ram[15041]  = 1;
  ram[15042]  = 1;
  ram[15043]  = 1;
  ram[15044]  = 1;
  ram[15045]  = 1;
  ram[15046]  = 1;
  ram[15047]  = 1;
  ram[15048]  = 1;
  ram[15049]  = 1;
  ram[15050]  = 1;
  ram[15051]  = 1;
  ram[15052]  = 1;
  ram[15053]  = 1;
  ram[15054]  = 1;
  ram[15055]  = 1;
  ram[15056]  = 1;
  ram[15057]  = 1;
  ram[15058]  = 1;
  ram[15059]  = 1;
  ram[15060]  = 1;
  ram[15061]  = 1;
  ram[15062]  = 1;
  ram[15063]  = 1;
  ram[15064]  = 1;
  ram[15065]  = 1;
  ram[15066]  = 1;
  ram[15067]  = 1;
  ram[15068]  = 1;
  ram[15069]  = 1;
  ram[15070]  = 1;
  ram[15071]  = 1;
  ram[15072]  = 1;
  ram[15073]  = 1;
  ram[15074]  = 1;
  ram[15075]  = 1;
  ram[15076]  = 1;
  ram[15077]  = 1;
  ram[15078]  = 1;
  ram[15079]  = 1;
  ram[15080]  = 1;
  ram[15081]  = 1;
  ram[15082]  = 1;
  ram[15083]  = 1;
  ram[15084]  = 1;
  ram[15085]  = 1;
  ram[15086]  = 1;
  ram[15087]  = 1;
  ram[15088]  = 1;
  ram[15089]  = 1;
  ram[15090]  = 1;
  ram[15091]  = 1;
  ram[15092]  = 1;
  ram[15093]  = 1;
  ram[15094]  = 1;
  ram[15095]  = 1;
  ram[15096]  = 1;
  ram[15097]  = 1;
  ram[15098]  = 1;
  ram[15099]  = 1;
  ram[15100]  = 1;
  ram[15101]  = 1;
  ram[15102]  = 1;
  ram[15103]  = 1;
  ram[15104]  = 1;
  ram[15105]  = 1;
  ram[15106]  = 1;
  ram[15107]  = 1;
  ram[15108]  = 1;
  ram[15109]  = 1;
  ram[15110]  = 1;
  ram[15111]  = 1;
  ram[15112]  = 1;
  ram[15113]  = 1;
  ram[15114]  = 1;
  ram[15115]  = 1;
  ram[15116]  = 1;
  ram[15117]  = 1;
  ram[15118]  = 1;
  ram[15119]  = 1;
  ram[15120]  = 1;
  ram[15121]  = 1;
  ram[15122]  = 1;
  ram[15123]  = 1;
  ram[15124]  = 1;
  ram[15125]  = 1;
  ram[15126]  = 1;
  ram[15127]  = 1;
  ram[15128]  = 1;
  ram[15129]  = 1;
  ram[15130]  = 1;
  ram[15131]  = 1;
  ram[15132]  = 1;
  ram[15133]  = 1;
  ram[15134]  = 1;
  ram[15135]  = 1;
  ram[15136]  = 1;
  ram[15137]  = 1;
  ram[15138]  = 1;
  ram[15139]  = 1;
  ram[15140]  = 1;
  ram[15141]  = 1;
  ram[15142]  = 1;
  ram[15143]  = 1;
  ram[15144]  = 1;
  ram[15145]  = 1;
  ram[15146]  = 1;
  ram[15147]  = 1;
  ram[15148]  = 1;
  ram[15149]  = 1;
  ram[15150]  = 1;
  ram[15151]  = 1;
  ram[15152]  = 1;
  ram[15153]  = 1;
  ram[15154]  = 1;
  ram[15155]  = 1;
  ram[15156]  = 1;
  ram[15157]  = 1;
  ram[15158]  = 1;
  ram[15159]  = 1;
  ram[15160]  = 1;
  ram[15161]  = 1;
  ram[15162]  = 1;
  ram[15163]  = 1;
  ram[15164]  = 1;
  ram[15165]  = 1;
  ram[15166]  = 1;
  ram[15167]  = 1;
  ram[15168]  = 1;
  ram[15169]  = 1;
  ram[15170]  = 1;
  ram[15171]  = 1;
  ram[15172]  = 1;
  ram[15173]  = 1;
  ram[15174]  = 1;
  ram[15175]  = 1;
  ram[15176]  = 1;
  ram[15177]  = 1;
  ram[15178]  = 1;
  ram[15179]  = 1;
  ram[15180]  = 1;
  ram[15181]  = 1;
  ram[15182]  = 1;
  ram[15183]  = 1;
  ram[15184]  = 1;
  ram[15185]  = 1;
  ram[15186]  = 1;
  ram[15187]  = 1;
  ram[15188]  = 1;
  ram[15189]  = 1;
  ram[15190]  = 1;
  ram[15191]  = 1;
  ram[15192]  = 1;
  ram[15193]  = 1;
  ram[15194]  = 1;
  ram[15195]  = 1;
  ram[15196]  = 1;
  ram[15197]  = 1;
  ram[15198]  = 1;
  ram[15199]  = 1;
  ram[15200]  = 1;
  ram[15201]  = 1;
  ram[15202]  = 1;
  ram[15203]  = 1;
  ram[15204]  = 1;
  ram[15205]  = 1;
  ram[15206]  = 1;
  ram[15207]  = 1;
  ram[15208]  = 1;
  ram[15209]  = 1;
  ram[15210]  = 1;
  ram[15211]  = 1;
  ram[15212]  = 1;
  ram[15213]  = 1;
  ram[15214]  = 1;
  ram[15215]  = 1;
  ram[15216]  = 1;
  ram[15217]  = 1;
  ram[15218]  = 1;
  ram[15219]  = 1;
  ram[15220]  = 1;
  ram[15221]  = 1;
  ram[15222]  = 1;
  ram[15223]  = 1;
  ram[15224]  = 1;
  ram[15225]  = 1;
  ram[15226]  = 1;
  ram[15227]  = 1;
  ram[15228]  = 1;
  ram[15229]  = 1;
  ram[15230]  = 1;
  ram[15231]  = 1;
  ram[15232]  = 1;
  ram[15233]  = 1;
  ram[15234]  = 1;
  ram[15235]  = 1;
  ram[15236]  = 1;
  ram[15237]  = 1;
  ram[15238]  = 1;
  ram[15239]  = 1;
  ram[15240]  = 1;
  ram[15241]  = 1;
  ram[15242]  = 1;
  ram[15243]  = 1;
  ram[15244]  = 1;
  ram[15245]  = 1;
  ram[15246]  = 1;
  ram[15247]  = 1;
  ram[15248]  = 1;
  ram[15249]  = 1;
  ram[15250]  = 1;
  ram[15251]  = 1;
  ram[15252]  = 1;
  ram[15253]  = 1;
  ram[15254]  = 1;
  ram[15255]  = 1;
  ram[15256]  = 1;
  ram[15257]  = 1;
  ram[15258]  = 1;
  ram[15259]  = 1;
  ram[15260]  = 1;
  ram[15261]  = 1;
  ram[15262]  = 1;
  ram[15263]  = 1;
  ram[15264]  = 1;
  ram[15265]  = 1;
  ram[15266]  = 1;
  ram[15267]  = 1;
  ram[15268]  = 1;
  ram[15269]  = 1;
  ram[15270]  = 1;
  ram[15271]  = 1;
  ram[15272]  = 1;
  ram[15273]  = 1;
  ram[15274]  = 1;
  ram[15275]  = 1;
  ram[15276]  = 1;
  ram[15277]  = 1;
  ram[15278]  = 1;
  ram[15279]  = 1;
  ram[15280]  = 1;
  ram[15281]  = 1;
  ram[15282]  = 1;
  ram[15283]  = 1;
  ram[15284]  = 1;
  ram[15285]  = 1;
  ram[15286]  = 1;
  ram[15287]  = 1;
  ram[15288]  = 1;
  ram[15289]  = 1;
  ram[15290]  = 1;
  ram[15291]  = 1;
  ram[15292]  = 1;
  ram[15293]  = 1;
  ram[15294]  = 1;
  ram[15295]  = 1;
  ram[15296]  = 1;
  ram[15297]  = 1;
  ram[15298]  = 1;
  ram[15299]  = 1;
  ram[15300]  = 1;
  ram[15301]  = 1;
  ram[15302]  = 1;
  ram[15303]  = 1;
  ram[15304]  = 1;
  ram[15305]  = 1;
  ram[15306]  = 1;
  ram[15307]  = 1;
  ram[15308]  = 1;
  ram[15309]  = 1;
  ram[15310]  = 1;
  ram[15311]  = 1;
  ram[15312]  = 1;
  ram[15313]  = 1;
  ram[15314]  = 1;
  ram[15315]  = 1;
  ram[15316]  = 1;
  ram[15317]  = 1;
  ram[15318]  = 1;
  ram[15319]  = 1;
  ram[15320]  = 1;
  ram[15321]  = 1;
  ram[15322]  = 1;
  ram[15323]  = 1;
  ram[15324]  = 1;
  ram[15325]  = 1;
  ram[15326]  = 1;
  ram[15327]  = 1;
  ram[15328]  = 1;
  ram[15329]  = 1;
  ram[15330]  = 1;
  ram[15331]  = 1;
  ram[15332]  = 1;
  ram[15333]  = 1;
  ram[15334]  = 1;
  ram[15335]  = 1;
  ram[15336]  = 1;
  ram[15337]  = 1;
  ram[15338]  = 1;
  ram[15339]  = 1;
  ram[15340]  = 1;
  ram[15341]  = 1;
  ram[15342]  = 1;
  ram[15343]  = 1;
  ram[15344]  = 1;
  ram[15345]  = 1;
  ram[15346]  = 1;
  ram[15347]  = 1;
  ram[15348]  = 1;
  ram[15349]  = 1;
  ram[15350]  = 1;
  ram[15351]  = 1;
  ram[15352]  = 1;
  ram[15353]  = 1;
  ram[15354]  = 1;
  ram[15355]  = 1;
  ram[15356]  = 1;
  ram[15357]  = 1;
  ram[15358]  = 1;
  ram[15359]  = 1;
  ram[15360]  = 1;
  ram[15361]  = 1;
  ram[15362]  = 1;
  ram[15363]  = 1;
  ram[15364]  = 1;
  ram[15365]  = 1;
  ram[15366]  = 1;
  ram[15367]  = 1;
  ram[15368]  = 1;
  ram[15369]  = 1;
  ram[15370]  = 1;
  ram[15371]  = 1;
  ram[15372]  = 1;
  ram[15373]  = 1;
  ram[15374]  = 1;
  ram[15375]  = 1;
  ram[15376]  = 1;
  ram[15377]  = 1;
  ram[15378]  = 1;
  ram[15379]  = 1;
  ram[15380]  = 1;
  ram[15381]  = 1;
  ram[15382]  = 1;
  ram[15383]  = 1;
  ram[15384]  = 1;
  ram[15385]  = 1;
  ram[15386]  = 1;
  ram[15387]  = 1;
  ram[15388]  = 1;
  ram[15389]  = 1;
  ram[15390]  = 1;
  ram[15391]  = 1;
  ram[15392]  = 1;
  ram[15393]  = 1;
  ram[15394]  = 1;
  ram[15395]  = 1;
  ram[15396]  = 1;
  ram[15397]  = 1;
  ram[15398]  = 1;
  ram[15399]  = 1;
  ram[15400]  = 1;
  ram[15401]  = 1;
  ram[15402]  = 1;
  ram[15403]  = 1;
  ram[15404]  = 1;
  ram[15405]  = 1;
  ram[15406]  = 1;
  ram[15407]  = 1;
  ram[15408]  = 1;
  ram[15409]  = 1;
  ram[15410]  = 1;
  ram[15411]  = 1;
  ram[15412]  = 1;
  ram[15413]  = 1;
  ram[15414]  = 1;
  ram[15415]  = 1;
  ram[15416]  = 1;
  ram[15417]  = 1;
  ram[15418]  = 1;
  ram[15419]  = 1;
  ram[15420]  = 1;
  ram[15421]  = 1;
  ram[15422]  = 1;
  ram[15423]  = 1;
  ram[15424]  = 1;
  ram[15425]  = 1;
  ram[15426]  = 1;
  ram[15427]  = 1;
  ram[15428]  = 1;
  ram[15429]  = 1;
  ram[15430]  = 1;
  ram[15431]  = 1;
  ram[15432]  = 1;
  ram[15433]  = 1;
  ram[15434]  = 1;
  ram[15435]  = 1;
  ram[15436]  = 1;
  ram[15437]  = 1;
  ram[15438]  = 1;
  ram[15439]  = 1;
  ram[15440]  = 1;
  ram[15441]  = 1;
  ram[15442]  = 1;
  ram[15443]  = 1;
  ram[15444]  = 1;
  ram[15445]  = 1;
  ram[15446]  = 1;
  ram[15447]  = 1;
  ram[15448]  = 1;
  ram[15449]  = 1;
  ram[15450]  = 1;
  ram[15451]  = 1;
  ram[15452]  = 1;
  ram[15453]  = 1;
  ram[15454]  = 1;
  ram[15455]  = 1;
  ram[15456]  = 1;
  ram[15457]  = 1;
  ram[15458]  = 1;
  ram[15459]  = 1;
  ram[15460]  = 1;
  ram[15461]  = 1;
  ram[15462]  = 1;
  ram[15463]  = 1;
  ram[15464]  = 1;
  ram[15465]  = 1;
  ram[15466]  = 1;
  ram[15467]  = 1;
  ram[15468]  = 1;
  ram[15469]  = 1;
  ram[15470]  = 1;
  ram[15471]  = 1;
  ram[15472]  = 1;
  ram[15473]  = 1;
  ram[15474]  = 1;
  ram[15475]  = 1;
  ram[15476]  = 1;
  ram[15477]  = 1;
  ram[15478]  = 1;
  ram[15479]  = 1;
  ram[15480]  = 1;
  ram[15481]  = 1;
  ram[15482]  = 1;
  ram[15483]  = 1;
  ram[15484]  = 1;
  ram[15485]  = 1;
  ram[15486]  = 1;
  ram[15487]  = 1;
  ram[15488]  = 1;
  ram[15489]  = 1;
  ram[15490]  = 1;
  ram[15491]  = 1;
  ram[15492]  = 1;
  ram[15493]  = 1;
  ram[15494]  = 1;
  ram[15495]  = 1;
  ram[15496]  = 1;
  ram[15497]  = 1;
  ram[15498]  = 1;
  ram[15499]  = 1;
  ram[15500]  = 1;
  ram[15501]  = 1;
  ram[15502]  = 1;
  ram[15503]  = 1;
  ram[15504]  = 1;
  ram[15505]  = 1;
  ram[15506]  = 1;
  ram[15507]  = 1;
  ram[15508]  = 1;
  ram[15509]  = 1;
  ram[15510]  = 1;
  ram[15511]  = 1;
  ram[15512]  = 1;
  ram[15513]  = 1;
  ram[15514]  = 1;
  ram[15515]  = 1;
  ram[15516]  = 1;
  ram[15517]  = 1;
  ram[15518]  = 1;
  ram[15519]  = 1;
  ram[15520]  = 1;
  ram[15521]  = 1;
  ram[15522]  = 1;
  ram[15523]  = 1;
  ram[15524]  = 1;
  ram[15525]  = 1;
  ram[15526]  = 1;
  ram[15527]  = 1;
  ram[15528]  = 1;
  ram[15529]  = 1;
  ram[15530]  = 1;
  ram[15531]  = 1;
  ram[15532]  = 1;
  ram[15533]  = 1;
  ram[15534]  = 1;
  ram[15535]  = 1;
  ram[15536]  = 1;
  ram[15537]  = 1;
  ram[15538]  = 1;
  ram[15539]  = 1;
  ram[15540]  = 1;
  ram[15541]  = 1;
  ram[15542]  = 1;
  ram[15543]  = 1;
  ram[15544]  = 1;
  ram[15545]  = 1;
  ram[15546]  = 1;
  ram[15547]  = 1;
  ram[15548]  = 1;
  ram[15549]  = 1;
  ram[15550]  = 1;
  ram[15551]  = 1;
  ram[15552]  = 1;
  ram[15553]  = 1;
  ram[15554]  = 1;
  ram[15555]  = 1;
  ram[15556]  = 1;
  ram[15557]  = 1;
  ram[15558]  = 1;
  ram[15559]  = 1;
  ram[15560]  = 1;
  ram[15561]  = 1;
  ram[15562]  = 1;
  ram[15563]  = 1;
  ram[15564]  = 1;
  ram[15565]  = 1;
  ram[15566]  = 1;
  ram[15567]  = 1;
  ram[15568]  = 1;
  ram[15569]  = 1;
  ram[15570]  = 1;
  ram[15571]  = 1;
  ram[15572]  = 1;
  ram[15573]  = 1;
  ram[15574]  = 1;
  ram[15575]  = 1;
  ram[15576]  = 1;
  ram[15577]  = 1;
  ram[15578]  = 1;
  ram[15579]  = 1;
  ram[15580]  = 1;
  ram[15581]  = 1;
  ram[15582]  = 1;
  ram[15583]  = 1;
  ram[15584]  = 1;
  ram[15585]  = 1;
  ram[15586]  = 1;
  ram[15587]  = 1;
  ram[15588]  = 1;
  ram[15589]  = 1;
  ram[15590]  = 1;
  ram[15591]  = 1;
  ram[15592]  = 1;
  ram[15593]  = 1;
  ram[15594]  = 1;
  ram[15595]  = 1;
  ram[15596]  = 1;
  ram[15597]  = 1;
  ram[15598]  = 1;
  ram[15599]  = 1;
  ram[15600]  = 1;
  ram[15601]  = 1;
  ram[15602]  = 1;
  ram[15603]  = 1;
  ram[15604]  = 1;
  ram[15605]  = 1;
  ram[15606]  = 1;
  ram[15607]  = 1;
  ram[15608]  = 1;
  ram[15609]  = 1;
  ram[15610]  = 1;
  ram[15611]  = 1;
  ram[15612]  = 1;
  ram[15613]  = 1;
  ram[15614]  = 1;
  ram[15615]  = 1;
  ram[15616]  = 1;
  ram[15617]  = 1;
  ram[15618]  = 1;
  ram[15619]  = 1;
  ram[15620]  = 1;
  ram[15621]  = 1;
  ram[15622]  = 1;
  ram[15623]  = 1;
  ram[15624]  = 1;
  ram[15625]  = 1;
  ram[15626]  = 1;
  ram[15627]  = 1;
  ram[15628]  = 1;
  ram[15629]  = 1;
  ram[15630]  = 1;
  ram[15631]  = 1;
  ram[15632]  = 1;
  ram[15633]  = 1;
  ram[15634]  = 1;
  ram[15635]  = 1;
  ram[15636]  = 1;
  ram[15637]  = 1;
  ram[15638]  = 1;
  ram[15639]  = 1;
  ram[15640]  = 1;
  ram[15641]  = 1;
  ram[15642]  = 1;
  ram[15643]  = 1;
  ram[15644]  = 1;
  ram[15645]  = 1;
  ram[15646]  = 1;
  ram[15647]  = 1;
  ram[15648]  = 1;
  ram[15649]  = 1;
  ram[15650]  = 1;
  ram[15651]  = 1;
  ram[15652]  = 1;
  ram[15653]  = 1;
  ram[15654]  = 1;
  ram[15655]  = 1;
  ram[15656]  = 1;
  ram[15657]  = 1;
  ram[15658]  = 1;
  ram[15659]  = 1;
  ram[15660]  = 1;
  ram[15661]  = 1;
  ram[15662]  = 1;
  ram[15663]  = 1;
  ram[15664]  = 1;
  ram[15665]  = 1;
  ram[15666]  = 1;
  ram[15667]  = 1;
  ram[15668]  = 1;
  ram[15669]  = 1;
  ram[15670]  = 1;
  ram[15671]  = 1;
  ram[15672]  = 1;
  ram[15673]  = 1;
  ram[15674]  = 1;
  ram[15675]  = 1;
  ram[15676]  = 1;
  ram[15677]  = 1;
  ram[15678]  = 1;
  ram[15679]  = 1;
  ram[15680]  = 1;
  ram[15681]  = 1;
  ram[15682]  = 1;
  ram[15683]  = 1;
  ram[15684]  = 1;
  ram[15685]  = 1;
  ram[15686]  = 1;
  ram[15687]  = 1;
  ram[15688]  = 1;
  ram[15689]  = 1;
  ram[15690]  = 1;
  ram[15691]  = 1;
  ram[15692]  = 1;
  ram[15693]  = 1;
  ram[15694]  = 1;
  ram[15695]  = 1;
  ram[15696]  = 1;
  ram[15697]  = 1;
  ram[15698]  = 1;
  ram[15699]  = 1;
  ram[15700]  = 1;
  ram[15701]  = 1;
  ram[15702]  = 1;
  ram[15703]  = 1;
  ram[15704]  = 1;
  ram[15705]  = 1;
  ram[15706]  = 1;
  ram[15707]  = 1;
  ram[15708]  = 1;
  ram[15709]  = 1;
  ram[15710]  = 1;
  ram[15711]  = 1;
  ram[15712]  = 1;
  ram[15713]  = 1;
  ram[15714]  = 1;
  ram[15715]  = 1;
  ram[15716]  = 1;
  ram[15717]  = 1;
  ram[15718]  = 1;
  ram[15719]  = 1;
  ram[15720]  = 1;
  ram[15721]  = 1;
  ram[15722]  = 1;
  ram[15723]  = 1;
  ram[15724]  = 1;
  ram[15725]  = 1;
  ram[15726]  = 1;
  ram[15727]  = 1;
  ram[15728]  = 1;
  ram[15729]  = 1;
  ram[15730]  = 1;
  ram[15731]  = 1;
  ram[15732]  = 1;
  ram[15733]  = 1;
  ram[15734]  = 1;
  ram[15735]  = 1;
  ram[15736]  = 1;
  ram[15737]  = 1;
  ram[15738]  = 1;
  ram[15739]  = 1;
  ram[15740]  = 1;
  ram[15741]  = 1;
  ram[15742]  = 1;
  ram[15743]  = 1;
  ram[15744]  = 1;
  ram[15745]  = 1;
  ram[15746]  = 1;
  ram[15747]  = 1;
  ram[15748]  = 1;
  ram[15749]  = 1;
  ram[15750]  = 1;
  ram[15751]  = 1;
  ram[15752]  = 1;
  ram[15753]  = 1;
  ram[15754]  = 1;
  ram[15755]  = 1;
  ram[15756]  = 1;
  ram[15757]  = 1;
  ram[15758]  = 1;
  ram[15759]  = 1;
  ram[15760]  = 1;
  ram[15761]  = 1;
  ram[15762]  = 1;
  ram[15763]  = 1;
  ram[15764]  = 1;
  ram[15765]  = 1;
  ram[15766]  = 1;
  ram[15767]  = 1;
  ram[15768]  = 1;
  ram[15769]  = 1;
  ram[15770]  = 1;
  ram[15771]  = 1;
  ram[15772]  = 1;
  ram[15773]  = 1;
  ram[15774]  = 1;
  ram[15775]  = 1;
  ram[15776]  = 1;
  ram[15777]  = 1;
  ram[15778]  = 1;
  ram[15779]  = 1;
  ram[15780]  = 1;
  ram[15781]  = 1;
  ram[15782]  = 1;
  ram[15783]  = 1;
  ram[15784]  = 1;
  ram[15785]  = 1;
  ram[15786]  = 1;
  ram[15787]  = 1;
  ram[15788]  = 1;
  ram[15789]  = 1;
  ram[15790]  = 1;
  ram[15791]  = 1;
  ram[15792]  = 1;
  ram[15793]  = 1;
  ram[15794]  = 1;
  ram[15795]  = 1;
  ram[15796]  = 1;
  ram[15797]  = 1;
  ram[15798]  = 1;
  ram[15799]  = 1;
  ram[15800]  = 1;
  ram[15801]  = 1;
  ram[15802]  = 1;
  ram[15803]  = 1;
  ram[15804]  = 1;
  ram[15805]  = 1;
  ram[15806]  = 1;
  ram[15807]  = 1;
  ram[15808]  = 1;
  ram[15809]  = 1;
  ram[15810]  = 1;
  ram[15811]  = 1;
  ram[15812]  = 1;
  ram[15813]  = 1;
  ram[15814]  = 1;
  ram[15815]  = 1;
  ram[15816]  = 1;
  ram[15817]  = 1;
  ram[15818]  = 1;
  ram[15819]  = 1;
  ram[15820]  = 1;
  ram[15821]  = 1;
  ram[15822]  = 1;
  ram[15823]  = 1;
  ram[15824]  = 1;
  ram[15825]  = 1;
  ram[15826]  = 1;
  ram[15827]  = 1;
  ram[15828]  = 1;
  ram[15829]  = 1;
  ram[15830]  = 1;
  ram[15831]  = 1;
  ram[15832]  = 1;
  ram[15833]  = 1;
  ram[15834]  = 1;
  ram[15835]  = 1;
  ram[15836]  = 1;
  ram[15837]  = 1;
  ram[15838]  = 1;
  ram[15839]  = 1;
  ram[15840]  = 1;
  ram[15841]  = 1;
  ram[15842]  = 1;
  ram[15843]  = 1;
  ram[15844]  = 1;
  ram[15845]  = 1;
  ram[15846]  = 1;
  ram[15847]  = 1;
  ram[15848]  = 1;
  ram[15849]  = 1;
  ram[15850]  = 1;
  ram[15851]  = 1;
  ram[15852]  = 1;
  ram[15853]  = 1;
  ram[15854]  = 1;
  ram[15855]  = 1;
  ram[15856]  = 1;
  ram[15857]  = 1;
  ram[15858]  = 1;
  ram[15859]  = 1;
  ram[15860]  = 1;
  ram[15861]  = 1;
  ram[15862]  = 1;
  ram[15863]  = 1;
  ram[15864]  = 1;
  ram[15865]  = 1;
  ram[15866]  = 1;
  ram[15867]  = 1;
  ram[15868]  = 1;
  ram[15869]  = 1;
  ram[15870]  = 1;
  ram[15871]  = 1;
  ram[15872]  = 1;
  ram[15873]  = 1;
  ram[15874]  = 1;
  ram[15875]  = 1;
  ram[15876]  = 1;
  ram[15877]  = 1;
  ram[15878]  = 1;
  ram[15879]  = 1;
  ram[15880]  = 1;
  ram[15881]  = 1;
  ram[15882]  = 1;
  ram[15883]  = 1;
  ram[15884]  = 1;
  ram[15885]  = 1;
  ram[15886]  = 1;
  ram[15887]  = 1;
  ram[15888]  = 1;
  ram[15889]  = 1;
  ram[15890]  = 1;
  ram[15891]  = 1;
  ram[15892]  = 1;
  ram[15893]  = 1;
  ram[15894]  = 1;
  ram[15895]  = 1;
  ram[15896]  = 1;
  ram[15897]  = 1;
  ram[15898]  = 1;
  ram[15899]  = 1;
  ram[15900]  = 1;
  ram[15901]  = 1;
  ram[15902]  = 1;
  ram[15903]  = 1;
  ram[15904]  = 1;
  ram[15905]  = 1;
  ram[15906]  = 1;
  ram[15907]  = 1;
  ram[15908]  = 1;
  ram[15909]  = 1;
  ram[15910]  = 1;
  ram[15911]  = 1;
  ram[15912]  = 1;
  ram[15913]  = 1;
  ram[15914]  = 1;
  ram[15915]  = 1;
  ram[15916]  = 1;
  ram[15917]  = 1;
  ram[15918]  = 1;
  ram[15919]  = 1;
  ram[15920]  = 1;
  ram[15921]  = 1;
  ram[15922]  = 1;
  ram[15923]  = 1;
  ram[15924]  = 1;
  ram[15925]  = 1;
  ram[15926]  = 1;
  ram[15927]  = 1;
  ram[15928]  = 1;
  ram[15929]  = 1;
  ram[15930]  = 1;
  ram[15931]  = 1;
  ram[15932]  = 1;
  ram[15933]  = 1;
  ram[15934]  = 1;
  ram[15935]  = 1;
  ram[15936]  = 1;
  ram[15937]  = 1;
  ram[15938]  = 1;
  ram[15939]  = 1;
  ram[15940]  = 1;
  ram[15941]  = 1;
  ram[15942]  = 1;
  ram[15943]  = 1;
  ram[15944]  = 1;
  ram[15945]  = 1;
  ram[15946]  = 1;
  ram[15947]  = 1;
  ram[15948]  = 1;
  ram[15949]  = 1;
  ram[15950]  = 1;
  ram[15951]  = 1;
  ram[15952]  = 1;
  ram[15953]  = 1;
  ram[15954]  = 1;
  ram[15955]  = 1;
  ram[15956]  = 1;
  ram[15957]  = 1;
  ram[15958]  = 1;
  ram[15959]  = 1;
  ram[15960]  = 1;
  ram[15961]  = 1;
  ram[15962]  = 1;
  ram[15963]  = 1;
  ram[15964]  = 1;
  ram[15965]  = 1;
  ram[15966]  = 1;
  ram[15967]  = 1;
  ram[15968]  = 1;
  ram[15969]  = 1;
  ram[15970]  = 1;
  ram[15971]  = 1;
  ram[15972]  = 1;
  ram[15973]  = 1;
  ram[15974]  = 1;
  ram[15975]  = 1;
  ram[15976]  = 1;
  ram[15977]  = 1;
  ram[15978]  = 1;
  ram[15979]  = 1;
  ram[15980]  = 1;
  ram[15981]  = 1;
  ram[15982]  = 1;
  ram[15983]  = 1;
  ram[15984]  = 1;
  ram[15985]  = 1;
  ram[15986]  = 1;
  ram[15987]  = 1;
  ram[15988]  = 1;
  ram[15989]  = 1;
  ram[15990]  = 1;
  ram[15991]  = 1;
  ram[15992]  = 1;
  ram[15993]  = 1;
  ram[15994]  = 1;
  ram[15995]  = 1;
  ram[15996]  = 1;
  ram[15997]  = 1;
  ram[15998]  = 1;
  ram[15999]  = 1;
  ram[16000]  = 1;
  ram[16001]  = 1;
  ram[16002]  = 1;
  ram[16003]  = 1;
  ram[16004]  = 1;
  ram[16005]  = 1;
  ram[16006]  = 1;
  ram[16007]  = 1;
  ram[16008]  = 1;
  ram[16009]  = 1;
  ram[16010]  = 1;
  ram[16011]  = 1;
  ram[16012]  = 1;
  ram[16013]  = 1;
  ram[16014]  = 1;
  ram[16015]  = 1;
  ram[16016]  = 1;
  ram[16017]  = 1;
  ram[16018]  = 1;
  ram[16019]  = 1;
  ram[16020]  = 1;
  ram[16021]  = 1;
  ram[16022]  = 1;
  ram[16023]  = 1;
  ram[16024]  = 1;
  ram[16025]  = 1;
  ram[16026]  = 1;
  ram[16027]  = 1;
  ram[16028]  = 1;
  ram[16029]  = 1;
  ram[16030]  = 1;
  ram[16031]  = 1;
  ram[16032]  = 1;
  ram[16033]  = 1;
  ram[16034]  = 1;
  ram[16035]  = 1;
  ram[16036]  = 1;
  ram[16037]  = 1;
  ram[16038]  = 1;
  ram[16039]  = 1;
  ram[16040]  = 1;
  ram[16041]  = 1;
  ram[16042]  = 1;
  ram[16043]  = 1;
  ram[16044]  = 1;
  ram[16045]  = 1;
  ram[16046]  = 1;
  ram[16047]  = 1;
  ram[16048]  = 1;
  ram[16049]  = 1;
  ram[16050]  = 1;
  ram[16051]  = 1;
  ram[16052]  = 1;
  ram[16053]  = 1;
  ram[16054]  = 1;
  ram[16055]  = 1;
  ram[16056]  = 1;
  ram[16057]  = 1;
  ram[16058]  = 1;
  ram[16059]  = 1;
  ram[16060]  = 1;
  ram[16061]  = 1;
  ram[16062]  = 1;
  ram[16063]  = 1;
  ram[16064]  = 1;
  ram[16065]  = 1;
  ram[16066]  = 1;
  ram[16067]  = 1;
  ram[16068]  = 1;
  ram[16069]  = 1;
  ram[16070]  = 1;
  ram[16071]  = 1;
  ram[16072]  = 1;
  ram[16073]  = 1;
  ram[16074]  = 1;
  ram[16075]  = 1;
  ram[16076]  = 1;
  ram[16077]  = 1;
  ram[16078]  = 1;
  ram[16079]  = 1;
  ram[16080]  = 1;
  ram[16081]  = 1;
  ram[16082]  = 1;
  ram[16083]  = 1;
  ram[16084]  = 1;
  ram[16085]  = 1;
  ram[16086]  = 1;
  ram[16087]  = 1;
  ram[16088]  = 1;
  ram[16089]  = 1;
  ram[16090]  = 1;
  ram[16091]  = 1;
  ram[16092]  = 1;
  ram[16093]  = 1;
  ram[16094]  = 1;
  ram[16095]  = 1;
  ram[16096]  = 1;
  ram[16097]  = 1;
  ram[16098]  = 1;
  ram[16099]  = 1;
  ram[16100]  = 1;
  ram[16101]  = 1;
  ram[16102]  = 1;
  ram[16103]  = 1;
  ram[16104]  = 1;
  ram[16105]  = 1;
  ram[16106]  = 1;
  ram[16107]  = 1;
  ram[16108]  = 1;
  ram[16109]  = 1;
  ram[16110]  = 1;
  ram[16111]  = 1;
  ram[16112]  = 1;
  ram[16113]  = 1;
  ram[16114]  = 1;
  ram[16115]  = 1;
  ram[16116]  = 1;
  ram[16117]  = 1;
  ram[16118]  = 1;
  ram[16119]  = 1;
  ram[16120]  = 1;
  ram[16121]  = 1;
  ram[16122]  = 1;
  ram[16123]  = 1;
  ram[16124]  = 1;
  ram[16125]  = 1;
  ram[16126]  = 1;
  ram[16127]  = 1;
  ram[16128]  = 1;
  ram[16129]  = 1;
  ram[16130]  = 1;
  ram[16131]  = 1;
  ram[16132]  = 1;
  ram[16133]  = 1;
  ram[16134]  = 1;
  ram[16135]  = 1;
  ram[16136]  = 1;
  ram[16137]  = 1;
  ram[16138]  = 1;
  ram[16139]  = 1;
  ram[16140]  = 1;
  ram[16141]  = 1;
  ram[16142]  = 1;
  ram[16143]  = 1;
  ram[16144]  = 1;
  ram[16145]  = 1;
  ram[16146]  = 1;
  ram[16147]  = 1;
  ram[16148]  = 1;
  ram[16149]  = 1;
  ram[16150]  = 1;
  ram[16151]  = 1;
  ram[16152]  = 1;
  ram[16153]  = 1;
  ram[16154]  = 1;
  ram[16155]  = 1;
  ram[16156]  = 1;
  ram[16157]  = 1;
  ram[16158]  = 1;
  ram[16159]  = 1;
  ram[16160]  = 1;
  ram[16161]  = 1;
  ram[16162]  = 1;
  ram[16163]  = 1;
  ram[16164]  = 1;
  ram[16165]  = 1;
  ram[16166]  = 1;
  ram[16167]  = 1;
  ram[16168]  = 1;
  ram[16169]  = 1;
  ram[16170]  = 1;
  ram[16171]  = 1;
  ram[16172]  = 1;
  ram[16173]  = 1;
  ram[16174]  = 1;
  ram[16175]  = 1;
  ram[16176]  = 1;
  ram[16177]  = 1;
  ram[16178]  = 1;
  ram[16179]  = 1;
  ram[16180]  = 1;
  ram[16181]  = 1;
  ram[16182]  = 1;
  ram[16183]  = 1;
  ram[16184]  = 1;
  ram[16185]  = 1;
  ram[16186]  = 1;
  ram[16187]  = 1;
  ram[16188]  = 1;
  ram[16189]  = 1;
  ram[16190]  = 1;
  ram[16191]  = 1;
  ram[16192]  = 1;
  ram[16193]  = 1;
  ram[16194]  = 1;
  ram[16195]  = 1;
  ram[16196]  = 1;
  ram[16197]  = 1;
  ram[16198]  = 1;
  ram[16199]  = 1;
  ram[16200]  = 1;
  ram[16201]  = 1;
  ram[16202]  = 1;
  ram[16203]  = 1;
  ram[16204]  = 1;
  ram[16205]  = 1;
  ram[16206]  = 1;
  ram[16207]  = 1;
  ram[16208]  = 1;
  ram[16209]  = 1;
  ram[16210]  = 1;
  ram[16211]  = 1;
  ram[16212]  = 1;
  ram[16213]  = 1;
  ram[16214]  = 1;
  ram[16215]  = 1;
  ram[16216]  = 1;
  ram[16217]  = 1;
  ram[16218]  = 1;
  ram[16219]  = 1;
  ram[16220]  = 1;
  ram[16221]  = 1;
  ram[16222]  = 1;
  ram[16223]  = 1;
  ram[16224]  = 1;
  ram[16225]  = 1;
  ram[16226]  = 1;
  ram[16227]  = 1;
  ram[16228]  = 1;
  ram[16229]  = 1;
  ram[16230]  = 1;
  ram[16231]  = 1;
  ram[16232]  = 1;
  ram[16233]  = 1;
  ram[16234]  = 1;
  ram[16235]  = 1;
  ram[16236]  = 1;
  ram[16237]  = 1;
  ram[16238]  = 1;
  ram[16239]  = 1;
  ram[16240]  = 1;
  ram[16241]  = 1;
  ram[16242]  = 1;
  ram[16243]  = 1;
  ram[16244]  = 1;
  ram[16245]  = 1;
  ram[16246]  = 1;
  ram[16247]  = 1;
  ram[16248]  = 1;
  ram[16249]  = 1;
  ram[16250]  = 1;
  ram[16251]  = 1;
  ram[16252]  = 1;
  ram[16253]  = 1;
  ram[16254]  = 1;
  ram[16255]  = 1;
  ram[16256]  = 1;
  ram[16257]  = 1;
  ram[16258]  = 1;
  ram[16259]  = 1;
  ram[16260]  = 1;
  ram[16261]  = 1;
  ram[16262]  = 1;
  ram[16263]  = 1;
  ram[16264]  = 1;
  ram[16265]  = 1;
  ram[16266]  = 1;
  ram[16267]  = 1;
  ram[16268]  = 1;
  ram[16269]  = 1;
  ram[16270]  = 1;
  ram[16271]  = 1;
  ram[16272]  = 1;
  ram[16273]  = 1;
  ram[16274]  = 1;
  ram[16275]  = 1;
  ram[16276]  = 1;
  ram[16277]  = 1;
  ram[16278]  = 1;
  ram[16279]  = 1;
  ram[16280]  = 1;
  ram[16281]  = 1;
  ram[16282]  = 1;
  ram[16283]  = 1;
  ram[16284]  = 1;
  ram[16285]  = 1;
  ram[16286]  = 1;
  ram[16287]  = 1;
  ram[16288]  = 1;
  ram[16289]  = 1;
  ram[16290]  = 1;
  ram[16291]  = 1;
  ram[16292]  = 1;
  ram[16293]  = 1;
  ram[16294]  = 1;
  ram[16295]  = 1;
  ram[16296]  = 1;
  ram[16297]  = 1;
  ram[16298]  = 1;
  ram[16299]  = 1;
  ram[16300]  = 1;
  ram[16301]  = 1;
  ram[16302]  = 1;
  ram[16303]  = 1;
  ram[16304]  = 1;
  ram[16305]  = 1;
  ram[16306]  = 1;
  ram[16307]  = 1;
  ram[16308]  = 1;
  ram[16309]  = 1;
  ram[16310]  = 1;
  ram[16311]  = 1;
  ram[16312]  = 1;
  ram[16313]  = 1;
  ram[16314]  = 1;
  ram[16315]  = 1;
  ram[16316]  = 1;
  ram[16317]  = 1;
  ram[16318]  = 1;
  ram[16319]  = 1;
  ram[16320]  = 1;
  ram[16321]  = 1;
  ram[16322]  = 1;
  ram[16323]  = 1;
  ram[16324]  = 1;
  ram[16325]  = 1;
  ram[16326]  = 1;
  ram[16327]  = 1;
  ram[16328]  = 1;
  ram[16329]  = 1;
  ram[16330]  = 1;
  ram[16331]  = 1;
  ram[16332]  = 1;
  ram[16333]  = 1;
  ram[16334]  = 1;
  ram[16335]  = 1;
  ram[16336]  = 1;
  ram[16337]  = 1;
  ram[16338]  = 1;
  ram[16339]  = 1;
  ram[16340]  = 1;
  ram[16341]  = 1;
  ram[16342]  = 1;
  ram[16343]  = 1;
  ram[16344]  = 1;
  ram[16345]  = 1;
  ram[16346]  = 1;
  ram[16347]  = 1;
  ram[16348]  = 1;
  ram[16349]  = 1;
  ram[16350]  = 1;
  ram[16351]  = 1;
  ram[16352]  = 1;
  ram[16353]  = 1;
  ram[16354]  = 1;
  ram[16355]  = 1;
  ram[16356]  = 1;
  ram[16357]  = 1;
  ram[16358]  = 1;
  ram[16359]  = 1;
  ram[16360]  = 1;
  ram[16361]  = 1;
  ram[16362]  = 1;
  ram[16363]  = 1;
  ram[16364]  = 1;
  ram[16365]  = 1;
  ram[16366]  = 1;
  ram[16367]  = 1;
  ram[16368]  = 1;
  ram[16369]  = 1;
  ram[16370]  = 1;
  ram[16371]  = 1;
  ram[16372]  = 1;
  ram[16373]  = 1;
  ram[16374]  = 1;
  ram[16375]  = 1;
  ram[16376]  = 1;
  ram[16377]  = 1;
  ram[16378]  = 1;
  ram[16379]  = 1;
  ram[16380]  = 1;
  ram[16381]  = 1;
  ram[16382]  = 1;
  ram[16383]  = 1;
  ram[16384]  = 1;
  ram[16385]  = 1;
  ram[16386]  = 1;
  ram[16387]  = 1;
  ram[16388]  = 1;
  ram[16389]  = 1;
  ram[16390]  = 1;
  ram[16391]  = 1;
  ram[16392]  = 1;
  ram[16393]  = 1;
  ram[16394]  = 1;
  ram[16395]  = 1;
  ram[16396]  = 1;
  ram[16397]  = 1;
  ram[16398]  = 1;
  ram[16399]  = 1;
  ram[16400]  = 1;
  ram[16401]  = 1;
  ram[16402]  = 1;
  ram[16403]  = 1;
  ram[16404]  = 1;
  ram[16405]  = 1;
  ram[16406]  = 1;
  ram[16407]  = 1;
  ram[16408]  = 1;
  ram[16409]  = 1;
  ram[16410]  = 1;
  ram[16411]  = 1;
  ram[16412]  = 1;
  ram[16413]  = 1;
  ram[16414]  = 1;
  ram[16415]  = 1;
  ram[16416]  = 1;
  ram[16417]  = 1;
  ram[16418]  = 1;
  ram[16419]  = 1;
  ram[16420]  = 1;
  ram[16421]  = 1;
  ram[16422]  = 1;
  ram[16423]  = 1;
  ram[16424]  = 1;
  ram[16425]  = 1;
  ram[16426]  = 1;
  ram[16427]  = 1;
  ram[16428]  = 1;
  ram[16429]  = 1;
  ram[16430]  = 1;
  ram[16431]  = 1;
  ram[16432]  = 1;
  ram[16433]  = 1;
  ram[16434]  = 1;
  ram[16435]  = 1;
  ram[16436]  = 1;
  ram[16437]  = 1;
  ram[16438]  = 1;
  ram[16439]  = 1;
  ram[16440]  = 1;
  ram[16441]  = 1;
  ram[16442]  = 1;
  ram[16443]  = 1;
  ram[16444]  = 1;
  ram[16445]  = 1;
  ram[16446]  = 1;
  ram[16447]  = 1;
  ram[16448]  = 1;
  ram[16449]  = 1;
  ram[16450]  = 1;
  ram[16451]  = 1;
  ram[16452]  = 1;
  ram[16453]  = 1;
  ram[16454]  = 1;
  ram[16455]  = 1;
  ram[16456]  = 1;
  ram[16457]  = 1;
  ram[16458]  = 1;
  ram[16459]  = 1;
  ram[16460]  = 1;
  ram[16461]  = 1;
  ram[16462]  = 1;
  ram[16463]  = 1;
  ram[16464]  = 1;
  ram[16465]  = 1;
  ram[16466]  = 1;
  ram[16467]  = 1;
  ram[16468]  = 1;
  ram[16469]  = 1;
  ram[16470]  = 1;
  ram[16471]  = 1;
  ram[16472]  = 1;
  ram[16473]  = 1;
  ram[16474]  = 1;
  ram[16475]  = 1;
  ram[16476]  = 1;
  ram[16477]  = 1;
  ram[16478]  = 1;
  ram[16479]  = 1;
  ram[16480]  = 1;
  ram[16481]  = 1;
  ram[16482]  = 1;
  ram[16483]  = 1;
  ram[16484]  = 1;
  ram[16485]  = 1;
  ram[16486]  = 1;
  ram[16487]  = 1;
  ram[16488]  = 1;
  ram[16489]  = 1;
  ram[16490]  = 1;
  ram[16491]  = 1;
  ram[16492]  = 1;
  ram[16493]  = 1;
  ram[16494]  = 1;
  ram[16495]  = 1;
  ram[16496]  = 1;
  ram[16497]  = 1;
  ram[16498]  = 1;
  ram[16499]  = 1;
  ram[16500]  = 1;
  ram[16501]  = 1;
  ram[16502]  = 1;
  ram[16503]  = 1;
  ram[16504]  = 1;
  ram[16505]  = 1;
  ram[16506]  = 1;
  ram[16507]  = 1;
  ram[16508]  = 1;
  ram[16509]  = 1;
  ram[16510]  = 1;
  ram[16511]  = 1;
  ram[16512]  = 1;
  ram[16513]  = 1;
  ram[16514]  = 1;
  ram[16515]  = 1;
  ram[16516]  = 1;
  ram[16517]  = 1;
  ram[16518]  = 1;
  ram[16519]  = 1;
  ram[16520]  = 1;
  ram[16521]  = 1;
  ram[16522]  = 1;
  ram[16523]  = 1;
  ram[16524]  = 1;
  ram[16525]  = 1;
  ram[16526]  = 1;
  ram[16527]  = 1;
  ram[16528]  = 1;
  ram[16529]  = 1;
  ram[16530]  = 1;
  ram[16531]  = 1;
  ram[16532]  = 1;
  ram[16533]  = 1;
  ram[16534]  = 1;
  ram[16535]  = 1;
  ram[16536]  = 1;
  ram[16537]  = 1;
  ram[16538]  = 1;
  ram[16539]  = 1;
  ram[16540]  = 1;
  ram[16541]  = 1;
  ram[16542]  = 1;
  ram[16543]  = 1;
  ram[16544]  = 1;
  ram[16545]  = 1;
  ram[16546]  = 1;
  ram[16547]  = 1;
  ram[16548]  = 1;
  ram[16549]  = 1;
  ram[16550]  = 1;
  ram[16551]  = 1;
  ram[16552]  = 1;
  ram[16553]  = 1;
  ram[16554]  = 1;
  ram[16555]  = 1;
  ram[16556]  = 1;
  ram[16557]  = 1;
  ram[16558]  = 1;
  ram[16559]  = 1;
  ram[16560]  = 1;
  ram[16561]  = 1;
  ram[16562]  = 1;
  ram[16563]  = 1;
  ram[16564]  = 1;
  ram[16565]  = 1;
  ram[16566]  = 1;
  ram[16567]  = 1;
  ram[16568]  = 1;
  ram[16569]  = 1;
  ram[16570]  = 1;
  ram[16571]  = 1;
  ram[16572]  = 1;
  ram[16573]  = 1;
  ram[16574]  = 1;
  ram[16575]  = 1;
  ram[16576]  = 1;
  ram[16577]  = 1;
  ram[16578]  = 1;
  ram[16579]  = 1;
  ram[16580]  = 1;
  ram[16581]  = 1;
  ram[16582]  = 1;
  ram[16583]  = 1;
  ram[16584]  = 1;
  ram[16585]  = 1;
  ram[16586]  = 1;
  ram[16587]  = 1;
  ram[16588]  = 1;
  ram[16589]  = 1;
  ram[16590]  = 1;
  ram[16591]  = 1;
  ram[16592]  = 1;
  ram[16593]  = 1;
  ram[16594]  = 1;
  ram[16595]  = 1;
  ram[16596]  = 1;
  ram[16597]  = 1;
  ram[16598]  = 1;
  ram[16599]  = 1;
  ram[16600]  = 1;
  ram[16601]  = 1;
  ram[16602]  = 1;
  ram[16603]  = 1;
  ram[16604]  = 1;
  ram[16605]  = 1;
  ram[16606]  = 1;
  ram[16607]  = 1;
  ram[16608]  = 1;
  ram[16609]  = 1;
  ram[16610]  = 1;
  ram[16611]  = 1;
  ram[16612]  = 1;
  ram[16613]  = 1;
  ram[16614]  = 1;
  ram[16615]  = 1;
  ram[16616]  = 1;
  ram[16617]  = 1;
  ram[16618]  = 1;
  ram[16619]  = 1;
  ram[16620]  = 1;
  ram[16621]  = 1;
  ram[16622]  = 1;
  ram[16623]  = 1;
  ram[16624]  = 1;
  ram[16625]  = 1;
  ram[16626]  = 1;
  ram[16627]  = 1;
  ram[16628]  = 1;
  ram[16629]  = 1;
  ram[16630]  = 1;
  ram[16631]  = 1;
  ram[16632]  = 1;
  ram[16633]  = 1;
  ram[16634]  = 1;
  ram[16635]  = 1;
  ram[16636]  = 1;
  ram[16637]  = 1;
  ram[16638]  = 1;
  ram[16639]  = 1;
  ram[16640]  = 1;
  ram[16641]  = 1;
  ram[16642]  = 1;
  ram[16643]  = 1;
  ram[16644]  = 1;
  ram[16645]  = 1;
  ram[16646]  = 1;
  ram[16647]  = 1;
  ram[16648]  = 1;
  ram[16649]  = 1;
  ram[16650]  = 1;
  ram[16651]  = 1;
  ram[16652]  = 1;
  ram[16653]  = 1;
  ram[16654]  = 1;
  ram[16655]  = 1;
  ram[16656]  = 1;
  ram[16657]  = 1;
  ram[16658]  = 1;
  ram[16659]  = 1;
  ram[16660]  = 1;
  ram[16661]  = 1;
  ram[16662]  = 1;
  ram[16663]  = 1;
  ram[16664]  = 1;
  ram[16665]  = 1;
  ram[16666]  = 1;
  ram[16667]  = 1;
  ram[16668]  = 1;
  ram[16669]  = 1;
  ram[16670]  = 1;
  ram[16671]  = 1;
  ram[16672]  = 1;
  ram[16673]  = 1;
  ram[16674]  = 1;
  ram[16675]  = 1;
  ram[16676]  = 1;
  ram[16677]  = 1;
  ram[16678]  = 1;
  ram[16679]  = 1;
  ram[16680]  = 1;
  ram[16681]  = 1;
  ram[16682]  = 1;
  ram[16683]  = 1;
  ram[16684]  = 1;
  ram[16685]  = 1;
  ram[16686]  = 1;
  ram[16687]  = 1;
  ram[16688]  = 1;
  ram[16689]  = 1;
  ram[16690]  = 1;
  ram[16691]  = 1;
  ram[16692]  = 1;
  ram[16693]  = 1;
  ram[16694]  = 1;
  ram[16695]  = 1;
  ram[16696]  = 1;
  ram[16697]  = 1;
  ram[16698]  = 1;
  ram[16699]  = 1;
  ram[16700]  = 1;
  ram[16701]  = 1;
  ram[16702]  = 1;
  ram[16703]  = 1;
  ram[16704]  = 1;
  ram[16705]  = 1;
  ram[16706]  = 1;
  ram[16707]  = 1;
  ram[16708]  = 1;
  ram[16709]  = 1;
  ram[16710]  = 1;
  ram[16711]  = 1;
  ram[16712]  = 1;
  ram[16713]  = 1;
  ram[16714]  = 1;
  ram[16715]  = 1;
  ram[16716]  = 1;
  ram[16717]  = 1;
  ram[16718]  = 1;
  ram[16719]  = 1;
  ram[16720]  = 1;
  ram[16721]  = 1;
  ram[16722]  = 1;
  ram[16723]  = 1;
  ram[16724]  = 1;
  ram[16725]  = 1;
  ram[16726]  = 1;
  ram[16727]  = 1;
  ram[16728]  = 1;
  ram[16729]  = 1;
  ram[16730]  = 1;
  ram[16731]  = 1;
  ram[16732]  = 1;
  ram[16733]  = 1;
  ram[16734]  = 1;
  ram[16735]  = 1;
  ram[16736]  = 1;
  ram[16737]  = 1;
  ram[16738]  = 1;
  ram[16739]  = 1;
  ram[16740]  = 1;
  ram[16741]  = 1;
  ram[16742]  = 1;
  ram[16743]  = 1;
  ram[16744]  = 1;
  ram[16745]  = 1;
  ram[16746]  = 1;
  ram[16747]  = 1;
  ram[16748]  = 1;
  ram[16749]  = 1;
  ram[16750]  = 1;
  ram[16751]  = 1;
  ram[16752]  = 1;
  ram[16753]  = 1;
  ram[16754]  = 1;
  ram[16755]  = 1;
  ram[16756]  = 1;
  ram[16757]  = 1;
  ram[16758]  = 1;
  ram[16759]  = 1;
  ram[16760]  = 1;
  ram[16761]  = 1;
  ram[16762]  = 1;
  ram[16763]  = 1;
  ram[16764]  = 1;
  ram[16765]  = 1;
  ram[16766]  = 1;
  ram[16767]  = 1;
  ram[16768]  = 1;
  ram[16769]  = 1;
  ram[16770]  = 1;
  ram[16771]  = 1;
  ram[16772]  = 1;
  ram[16773]  = 1;
  ram[16774]  = 1;
  ram[16775]  = 1;
  ram[16776]  = 1;
  ram[16777]  = 1;
  ram[16778]  = 1;
  ram[16779]  = 1;
  ram[16780]  = 1;
  ram[16781]  = 1;
  ram[16782]  = 1;
  ram[16783]  = 1;
  ram[16784]  = 1;
  ram[16785]  = 1;
  ram[16786]  = 1;
  ram[16787]  = 1;
  ram[16788]  = 1;
  ram[16789]  = 1;
  ram[16790]  = 1;
  ram[16791]  = 1;
  ram[16792]  = 1;
  ram[16793]  = 1;
  ram[16794]  = 1;
  ram[16795]  = 1;
  ram[16796]  = 1;
  ram[16797]  = 1;
  ram[16798]  = 1;
  ram[16799]  = 1;
  ram[16800]  = 1;
  ram[16801]  = 1;
  ram[16802]  = 1;
  ram[16803]  = 1;
  ram[16804]  = 1;
  ram[16805]  = 1;
  ram[16806]  = 1;
  ram[16807]  = 1;
  ram[16808]  = 1;
  ram[16809]  = 1;
  ram[16810]  = 1;
  ram[16811]  = 1;
  ram[16812]  = 1;
  ram[16813]  = 1;
  ram[16814]  = 1;
  ram[16815]  = 1;
  ram[16816]  = 1;
  ram[16817]  = 1;
  ram[16818]  = 1;
  ram[16819]  = 1;
  ram[16820]  = 1;
  ram[16821]  = 1;
  ram[16822]  = 1;
  ram[16823]  = 1;
  ram[16824]  = 1;
  ram[16825]  = 1;
  ram[16826]  = 1;
  ram[16827]  = 1;
  ram[16828]  = 1;
  ram[16829]  = 1;
  ram[16830]  = 1;
  ram[16831]  = 1;
  ram[16832]  = 1;
  ram[16833]  = 1;
  ram[16834]  = 1;
  ram[16835]  = 1;
  ram[16836]  = 1;
  ram[16837]  = 1;
  ram[16838]  = 1;
  ram[16839]  = 1;
  ram[16840]  = 1;
  ram[16841]  = 1;
  ram[16842]  = 1;
  ram[16843]  = 1;
  ram[16844]  = 1;
  ram[16845]  = 1;
  ram[16846]  = 1;
  ram[16847]  = 1;
  ram[16848]  = 1;
  ram[16849]  = 1;
  ram[16850]  = 1;
  ram[16851]  = 1;
  ram[16852]  = 1;
  ram[16853]  = 1;
  ram[16854]  = 1;
  ram[16855]  = 1;
  ram[16856]  = 1;
  ram[16857]  = 1;
  ram[16858]  = 1;
  ram[16859]  = 1;
  ram[16860]  = 1;
  ram[16861]  = 1;
  ram[16862]  = 1;
  ram[16863]  = 1;
  ram[16864]  = 1;
  ram[16865]  = 1;
  ram[16866]  = 1;
  ram[16867]  = 1;
  ram[16868]  = 1;
  ram[16869]  = 1;
  ram[16870]  = 1;
  ram[16871]  = 1;
  ram[16872]  = 1;
  ram[16873]  = 1;
  ram[16874]  = 1;
  ram[16875]  = 1;
  ram[16876]  = 1;
  ram[16877]  = 1;
  ram[16878]  = 1;
  ram[16879]  = 1;
  ram[16880]  = 1;
  ram[16881]  = 1;
  ram[16882]  = 1;
  ram[16883]  = 1;
  ram[16884]  = 1;
  ram[16885]  = 1;
  ram[16886]  = 1;
  ram[16887]  = 1;
  ram[16888]  = 1;
  ram[16889]  = 1;
  ram[16890]  = 1;
  ram[16891]  = 1;
  ram[16892]  = 1;
  ram[16893]  = 1;
  ram[16894]  = 1;
  ram[16895]  = 1;
  ram[16896]  = 1;
  ram[16897]  = 1;
  ram[16898]  = 1;
  ram[16899]  = 1;
  ram[16900]  = 1;
  ram[16901]  = 1;
  ram[16902]  = 1;
  ram[16903]  = 1;
  ram[16904]  = 1;
  ram[16905]  = 1;
  ram[16906]  = 1;
  ram[16907]  = 1;
  ram[16908]  = 1;
  ram[16909]  = 1;
  ram[16910]  = 1;
  ram[16911]  = 1;
  ram[16912]  = 1;
  ram[16913]  = 1;
  ram[16914]  = 1;
  ram[16915]  = 1;
  ram[16916]  = 1;
  ram[16917]  = 1;
  ram[16918]  = 1;
  ram[16919]  = 1;
  ram[16920]  = 1;
  ram[16921]  = 1;
  ram[16922]  = 1;
  ram[16923]  = 1;
  ram[16924]  = 1;
  ram[16925]  = 1;
  ram[16926]  = 1;
  ram[16927]  = 1;
  ram[16928]  = 1;
  ram[16929]  = 1;
  ram[16930]  = 1;
  ram[16931]  = 1;
  ram[16932]  = 1;
  ram[16933]  = 1;
  ram[16934]  = 1;
  ram[16935]  = 1;
  ram[16936]  = 1;
  ram[16937]  = 1;
  ram[16938]  = 1;
  ram[16939]  = 1;
  ram[16940]  = 1;
  ram[16941]  = 1;
  ram[16942]  = 1;
  ram[16943]  = 1;
  ram[16944]  = 1;
  ram[16945]  = 1;
  ram[16946]  = 1;
  ram[16947]  = 1;
  ram[16948]  = 1;
  ram[16949]  = 1;
  ram[16950]  = 1;
  ram[16951]  = 1;
  ram[16952]  = 1;
  ram[16953]  = 1;
  ram[16954]  = 1;
  ram[16955]  = 1;
  ram[16956]  = 1;
  ram[16957]  = 1;
  ram[16958]  = 1;
  ram[16959]  = 1;
  ram[16960]  = 1;
  ram[16961]  = 1;
  ram[16962]  = 1;
  ram[16963]  = 1;
  ram[16964]  = 1;
  ram[16965]  = 1;
  ram[16966]  = 1;
  ram[16967]  = 1;
  ram[16968]  = 1;
  ram[16969]  = 1;
  ram[16970]  = 1;
  ram[16971]  = 1;
  ram[16972]  = 1;
  ram[16973]  = 1;
  ram[16974]  = 1;
  ram[16975]  = 1;
  ram[16976]  = 1;
  ram[16977]  = 1;
  ram[16978]  = 1;
  ram[16979]  = 1;
  ram[16980]  = 1;
  ram[16981]  = 1;
  ram[16982]  = 1;
  ram[16983]  = 1;
  ram[16984]  = 1;
  ram[16985]  = 1;
  ram[16986]  = 1;
  ram[16987]  = 1;
  ram[16988]  = 1;
  ram[16989]  = 1;
  ram[16990]  = 1;
  ram[16991]  = 1;
  ram[16992]  = 1;
  ram[16993]  = 1;
  ram[16994]  = 1;
  ram[16995]  = 1;
  ram[16996]  = 1;
  ram[16997]  = 1;
  ram[16998]  = 1;
  ram[16999]  = 1;
  ram[17000]  = 1;
  ram[17001]  = 1;
  ram[17002]  = 1;
  ram[17003]  = 1;
  ram[17004]  = 1;
  ram[17005]  = 1;
  ram[17006]  = 1;
  ram[17007]  = 1;
  ram[17008]  = 1;
  ram[17009]  = 1;
  ram[17010]  = 1;
  ram[17011]  = 1;
  ram[17012]  = 1;
  ram[17013]  = 1;
  ram[17014]  = 1;
  ram[17015]  = 1;
  ram[17016]  = 1;
  ram[17017]  = 1;
  ram[17018]  = 1;
  ram[17019]  = 1;
  ram[17020]  = 1;
  ram[17021]  = 1;
  ram[17022]  = 1;
  ram[17023]  = 1;
  ram[17024]  = 1;
  ram[17025]  = 1;
  ram[17026]  = 1;
  ram[17027]  = 1;
  ram[17028]  = 1;
  ram[17029]  = 1;
  ram[17030]  = 1;
  ram[17031]  = 1;
  ram[17032]  = 1;
  ram[17033]  = 1;
  ram[17034]  = 1;
  ram[17035]  = 1;
  ram[17036]  = 1;
  ram[17037]  = 1;
  ram[17038]  = 1;
  ram[17039]  = 1;
  ram[17040]  = 1;
  ram[17041]  = 1;
  ram[17042]  = 1;
  ram[17043]  = 1;
  ram[17044]  = 1;
  ram[17045]  = 1;
  ram[17046]  = 1;
  ram[17047]  = 1;
  ram[17048]  = 1;
  ram[17049]  = 1;
  ram[17050]  = 1;
  ram[17051]  = 1;
  ram[17052]  = 1;
  ram[17053]  = 1;
  ram[17054]  = 1;
  ram[17055]  = 1;
  ram[17056]  = 1;
  ram[17057]  = 1;
  ram[17058]  = 1;
  ram[17059]  = 1;
  ram[17060]  = 1;
  ram[17061]  = 1;
  ram[17062]  = 1;
  ram[17063]  = 1;
  ram[17064]  = 1;
  ram[17065]  = 1;
  ram[17066]  = 1;
  ram[17067]  = 1;
  ram[17068]  = 1;
  ram[17069]  = 1;
  ram[17070]  = 1;
  ram[17071]  = 1;
  ram[17072]  = 1;
  ram[17073]  = 1;
  ram[17074]  = 1;
  ram[17075]  = 1;
  ram[17076]  = 1;
  ram[17077]  = 1;
  ram[17078]  = 1;
  ram[17079]  = 1;
  ram[17080]  = 1;
  ram[17081]  = 1;
  ram[17082]  = 1;
  ram[17083]  = 1;
  ram[17084]  = 1;
  ram[17085]  = 1;
  ram[17086]  = 1;
  ram[17087]  = 1;
  ram[17088]  = 1;
  ram[17089]  = 1;
  ram[17090]  = 1;
  ram[17091]  = 1;
  ram[17092]  = 1;
  ram[17093]  = 1;
  ram[17094]  = 1;
  ram[17095]  = 1;
  ram[17096]  = 1;
  ram[17097]  = 1;
  ram[17098]  = 1;
  ram[17099]  = 1;
  ram[17100]  = 1;
  ram[17101]  = 1;
  ram[17102]  = 1;
  ram[17103]  = 1;
  ram[17104]  = 1;
  ram[17105]  = 1;
  ram[17106]  = 1;
  ram[17107]  = 1;
  ram[17108]  = 1;
  ram[17109]  = 1;
  ram[17110]  = 1;
  ram[17111]  = 1;
  ram[17112]  = 1;
  ram[17113]  = 1;
  ram[17114]  = 1;
  ram[17115]  = 1;
  ram[17116]  = 1;
  ram[17117]  = 1;
  ram[17118]  = 1;
  ram[17119]  = 1;
  ram[17120]  = 1;
  ram[17121]  = 1;
  ram[17122]  = 1;
  ram[17123]  = 1;
  ram[17124]  = 1;
  ram[17125]  = 1;
  ram[17126]  = 1;
  ram[17127]  = 1;
  ram[17128]  = 1;
  ram[17129]  = 1;
  ram[17130]  = 1;
  ram[17131]  = 1;
  ram[17132]  = 1;
  ram[17133]  = 1;
  ram[17134]  = 1;
  ram[17135]  = 1;
  ram[17136]  = 1;
  ram[17137]  = 1;
  ram[17138]  = 1;
  ram[17139]  = 1;
  ram[17140]  = 1;
  ram[17141]  = 1;
  ram[17142]  = 1;
  ram[17143]  = 1;
  ram[17144]  = 1;
  ram[17145]  = 1;
  ram[17146]  = 1;
  ram[17147]  = 1;
  ram[17148]  = 1;
  ram[17149]  = 1;
  ram[17150]  = 1;
  ram[17151]  = 1;
  ram[17152]  = 1;
  ram[17153]  = 1;
  ram[17154]  = 1;
  ram[17155]  = 1;
  ram[17156]  = 1;
  ram[17157]  = 1;
  ram[17158]  = 1;
  ram[17159]  = 1;
  ram[17160]  = 1;
  ram[17161]  = 1;
  ram[17162]  = 1;
  ram[17163]  = 1;
  ram[17164]  = 1;
  ram[17165]  = 1;
  ram[17166]  = 1;
  ram[17167]  = 1;
  ram[17168]  = 1;
  ram[17169]  = 1;
  ram[17170]  = 1;
  ram[17171]  = 1;
  ram[17172]  = 1;
  ram[17173]  = 1;
  ram[17174]  = 1;
  ram[17175]  = 1;
  ram[17176]  = 1;
  ram[17177]  = 1;
  ram[17178]  = 1;
  ram[17179]  = 1;
  ram[17180]  = 1;
  ram[17181]  = 1;
  ram[17182]  = 1;
  ram[17183]  = 1;
  ram[17184]  = 1;
  ram[17185]  = 1;
  ram[17186]  = 1;
  ram[17187]  = 1;
  ram[17188]  = 1;
  ram[17189]  = 1;
  ram[17190]  = 1;
  ram[17191]  = 1;
  ram[17192]  = 1;
  ram[17193]  = 1;
  ram[17194]  = 1;
  ram[17195]  = 1;
  ram[17196]  = 1;
  ram[17197]  = 1;
  ram[17198]  = 1;
  ram[17199]  = 1;
  ram[17200]  = 1;
  ram[17201]  = 1;
  ram[17202]  = 1;
  ram[17203]  = 1;
  ram[17204]  = 1;
  ram[17205]  = 1;
  ram[17206]  = 1;
  ram[17207]  = 1;
  ram[17208]  = 1;
  ram[17209]  = 1;
  ram[17210]  = 1;
  ram[17211]  = 1;
  ram[17212]  = 1;
  ram[17213]  = 1;
  ram[17214]  = 1;
  ram[17215]  = 1;
  ram[17216]  = 1;
  ram[17217]  = 1;
  ram[17218]  = 1;
  ram[17219]  = 1;
  ram[17220]  = 1;
  ram[17221]  = 1;
  ram[17222]  = 1;
  ram[17223]  = 1;
  ram[17224]  = 1;
  ram[17225]  = 1;
  ram[17226]  = 1;
  ram[17227]  = 1;
  ram[17228]  = 1;
  ram[17229]  = 1;
  ram[17230]  = 1;
  ram[17231]  = 1;
  ram[17232]  = 1;
  ram[17233]  = 1;
  ram[17234]  = 1;
  ram[17235]  = 1;
  ram[17236]  = 1;
  ram[17237]  = 1;
  ram[17238]  = 1;
  ram[17239]  = 1;
  ram[17240]  = 1;
  ram[17241]  = 1;
  ram[17242]  = 1;
  ram[17243]  = 1;
  ram[17244]  = 1;
  ram[17245]  = 1;
  ram[17246]  = 1;
  ram[17247]  = 1;
  ram[17248]  = 1;
  ram[17249]  = 1;
  ram[17250]  = 1;
  ram[17251]  = 1;
  ram[17252]  = 1;
  ram[17253]  = 1;
  ram[17254]  = 1;
  ram[17255]  = 1;
  ram[17256]  = 1;
  ram[17257]  = 1;
  ram[17258]  = 1;
  ram[17259]  = 1;
  ram[17260]  = 1;
  ram[17261]  = 1;
  ram[17262]  = 1;
  ram[17263]  = 1;
  ram[17264]  = 1;
  ram[17265]  = 1;
  ram[17266]  = 1;
  ram[17267]  = 1;
  ram[17268]  = 1;
  ram[17269]  = 1;
  ram[17270]  = 1;
  ram[17271]  = 1;
  ram[17272]  = 1;
  ram[17273]  = 1;
  ram[17274]  = 1;
  ram[17275]  = 1;
  ram[17276]  = 1;
  ram[17277]  = 1;
  ram[17278]  = 1;
  ram[17279]  = 1;
  ram[17280]  = 1;
  ram[17281]  = 1;
  ram[17282]  = 1;
  ram[17283]  = 1;
  ram[17284]  = 1;
  ram[17285]  = 1;
  ram[17286]  = 1;
  ram[17287]  = 1;
  ram[17288]  = 1;
  ram[17289]  = 1;
  ram[17290]  = 1;
  ram[17291]  = 1;
  ram[17292]  = 1;
  ram[17293]  = 1;
  ram[17294]  = 1;
  ram[17295]  = 1;
  ram[17296]  = 1;
  ram[17297]  = 1;
  ram[17298]  = 1;
  ram[17299]  = 1;
  ram[17300]  = 1;
  ram[17301]  = 1;
  ram[17302]  = 1;
  ram[17303]  = 1;
  ram[17304]  = 1;
  ram[17305]  = 1;
  ram[17306]  = 1;
  ram[17307]  = 1;
  ram[17308]  = 1;
  ram[17309]  = 1;
  ram[17310]  = 1;
  ram[17311]  = 1;
  ram[17312]  = 1;
  ram[17313]  = 1;
  ram[17314]  = 1;
  ram[17315]  = 1;
  ram[17316]  = 1;
  ram[17317]  = 1;
  ram[17318]  = 1;
  ram[17319]  = 1;
  ram[17320]  = 1;
  ram[17321]  = 1;
  ram[17322]  = 1;
  ram[17323]  = 1;
  ram[17324]  = 1;
  ram[17325]  = 1;
  ram[17326]  = 1;
  ram[17327]  = 1;
  ram[17328]  = 1;
  ram[17329]  = 1;
  ram[17330]  = 1;
  ram[17331]  = 1;
  ram[17332]  = 1;
  ram[17333]  = 1;
  ram[17334]  = 1;
  ram[17335]  = 1;
  ram[17336]  = 1;
  ram[17337]  = 1;
  ram[17338]  = 1;
  ram[17339]  = 1;
  ram[17340]  = 1;
  ram[17341]  = 1;
  ram[17342]  = 1;
  ram[17343]  = 1;
  ram[17344]  = 1;
  ram[17345]  = 1;
  ram[17346]  = 1;
  ram[17347]  = 1;
  ram[17348]  = 1;
  ram[17349]  = 1;
  ram[17350]  = 1;
  ram[17351]  = 1;
  ram[17352]  = 1;
  ram[17353]  = 1;
  ram[17354]  = 1;
  ram[17355]  = 1;
  ram[17356]  = 1;
  ram[17357]  = 1;
  ram[17358]  = 1;
  ram[17359]  = 1;
  ram[17360]  = 1;
  ram[17361]  = 1;
  ram[17362]  = 1;
  ram[17363]  = 1;
  ram[17364]  = 1;
  ram[17365]  = 1;
  ram[17366]  = 1;
  ram[17367]  = 1;
  ram[17368]  = 1;
  ram[17369]  = 1;
  ram[17370]  = 1;
  ram[17371]  = 1;
  ram[17372]  = 1;
  ram[17373]  = 1;
  ram[17374]  = 1;
  ram[17375]  = 1;
  ram[17376]  = 1;
  ram[17377]  = 1;
  ram[17378]  = 1;
  ram[17379]  = 1;
  ram[17380]  = 1;
  ram[17381]  = 1;
  ram[17382]  = 1;
  ram[17383]  = 1;
  ram[17384]  = 1;
  ram[17385]  = 1;
  ram[17386]  = 1;
  ram[17387]  = 1;
  ram[17388]  = 1;
  ram[17389]  = 1;
  ram[17390]  = 1;
  ram[17391]  = 1;
  ram[17392]  = 1;
  ram[17393]  = 1;
  ram[17394]  = 1;
  ram[17395]  = 1;
  ram[17396]  = 1;
  ram[17397]  = 1;
  ram[17398]  = 1;
  ram[17399]  = 1;
  ram[17400]  = 1;
  ram[17401]  = 1;
  ram[17402]  = 1;
  ram[17403]  = 1;
  ram[17404]  = 1;
  ram[17405]  = 1;
  ram[17406]  = 1;
  ram[17407]  = 1;
  ram[17408]  = 1;
  ram[17409]  = 1;
  ram[17410]  = 1;
  ram[17411]  = 1;
  ram[17412]  = 1;
  ram[17413]  = 1;
  ram[17414]  = 1;
  ram[17415]  = 1;
  ram[17416]  = 1;
  ram[17417]  = 1;
  ram[17418]  = 1;
  ram[17419]  = 1;
  ram[17420]  = 1;
  ram[17421]  = 1;
  ram[17422]  = 1;
  ram[17423]  = 1;
  ram[17424]  = 1;
  ram[17425]  = 1;
  ram[17426]  = 1;
  ram[17427]  = 1;
  ram[17428]  = 1;
  ram[17429]  = 1;
  ram[17430]  = 1;
  ram[17431]  = 1;
  ram[17432]  = 1;
  ram[17433]  = 1;
  ram[17434]  = 1;
  ram[17435]  = 1;
  ram[17436]  = 1;
  ram[17437]  = 1;
  ram[17438]  = 1;
  ram[17439]  = 1;
  ram[17440]  = 1;
  ram[17441]  = 1;
  ram[17442]  = 1;
  ram[17443]  = 1;
  ram[17444]  = 1;
  ram[17445]  = 1;
  ram[17446]  = 1;
  ram[17447]  = 1;
  ram[17448]  = 1;
  ram[17449]  = 1;
  ram[17450]  = 1;
  ram[17451]  = 1;
  ram[17452]  = 1;
  ram[17453]  = 1;
  ram[17454]  = 1;
  ram[17455]  = 1;
  ram[17456]  = 1;
  ram[17457]  = 1;
  ram[17458]  = 1;
  ram[17459]  = 1;
  ram[17460]  = 1;
  ram[17461]  = 1;
  ram[17462]  = 1;
  ram[17463]  = 1;
  ram[17464]  = 1;
  ram[17465]  = 1;
  ram[17466]  = 1;
  ram[17467]  = 1;
  ram[17468]  = 1;
  ram[17469]  = 1;
  ram[17470]  = 1;
  ram[17471]  = 1;
  ram[17472]  = 1;
  ram[17473]  = 1;
  ram[17474]  = 1;
  ram[17475]  = 1;
  ram[17476]  = 1;
  ram[17477]  = 1;
  ram[17478]  = 1;
  ram[17479]  = 1;
  ram[17480]  = 1;
  ram[17481]  = 1;
  ram[17482]  = 1;
  ram[17483]  = 1;
  ram[17484]  = 1;
  ram[17485]  = 1;
  ram[17486]  = 1;
  ram[17487]  = 1;
  ram[17488]  = 1;
  ram[17489]  = 1;
  ram[17490]  = 1;
  ram[17491]  = 1;
  ram[17492]  = 1;
  ram[17493]  = 1;
  ram[17494]  = 1;
  ram[17495]  = 1;
  ram[17496]  = 1;
  ram[17497]  = 1;
  ram[17498]  = 1;
  ram[17499]  = 1;
  ram[17500]  = 1;
  ram[17501]  = 1;
  ram[17502]  = 1;
  ram[17503]  = 1;
  ram[17504]  = 1;
  ram[17505]  = 1;
  ram[17506]  = 1;
  ram[17507]  = 1;
  ram[17508]  = 1;
  ram[17509]  = 1;
  ram[17510]  = 1;
  ram[17511]  = 1;
  ram[17512]  = 1;
  ram[17513]  = 1;
  ram[17514]  = 1;
  ram[17515]  = 1;
  ram[17516]  = 1;
  ram[17517]  = 1;
  ram[17518]  = 1;
  ram[17519]  = 1;
  ram[17520]  = 1;
  ram[17521]  = 1;
  ram[17522]  = 1;
  ram[17523]  = 1;
  ram[17524]  = 1;
  ram[17525]  = 1;
  ram[17526]  = 1;
  ram[17527]  = 1;
  ram[17528]  = 1;
  ram[17529]  = 1;
  ram[17530]  = 1;
  ram[17531]  = 1;
  ram[17532]  = 1;
  ram[17533]  = 1;
  ram[17534]  = 1;
  ram[17535]  = 1;
  ram[17536]  = 1;
  ram[17537]  = 1;
  ram[17538]  = 1;
  ram[17539]  = 1;
  ram[17540]  = 1;
  ram[17541]  = 1;
  ram[17542]  = 1;
  ram[17543]  = 1;
  ram[17544]  = 1;
  ram[17545]  = 1;
  ram[17546]  = 1;
  ram[17547]  = 1;
  ram[17548]  = 1;
  ram[17549]  = 1;
  ram[17550]  = 1;
  ram[17551]  = 1;
  ram[17552]  = 1;
  ram[17553]  = 1;
  ram[17554]  = 1;
  ram[17555]  = 1;
  ram[17556]  = 1;
  ram[17557]  = 1;
  ram[17558]  = 1;
  ram[17559]  = 1;
  ram[17560]  = 1;
  ram[17561]  = 1;
  ram[17562]  = 1;
  ram[17563]  = 1;
  ram[17564]  = 1;
  ram[17565]  = 1;
  ram[17566]  = 1;
  ram[17567]  = 1;
  ram[17568]  = 1;
  ram[17569]  = 1;
  ram[17570]  = 1;
  ram[17571]  = 1;
  ram[17572]  = 1;
  ram[17573]  = 1;
  ram[17574]  = 1;
  ram[17575]  = 1;
  ram[17576]  = 1;
  ram[17577]  = 1;
  ram[17578]  = 1;
  ram[17579]  = 1;
  ram[17580]  = 1;
  ram[17581]  = 1;
  ram[17582]  = 1;
  ram[17583]  = 1;
  ram[17584]  = 1;
  ram[17585]  = 1;
  ram[17586]  = 1;
  ram[17587]  = 1;
  ram[17588]  = 1;
  ram[17589]  = 1;
  ram[17590]  = 1;
  ram[17591]  = 1;
  ram[17592]  = 1;
  ram[17593]  = 1;
  ram[17594]  = 1;
  ram[17595]  = 1;
  ram[17596]  = 1;
  ram[17597]  = 1;
  ram[17598]  = 1;
  ram[17599]  = 1;
  ram[17600]  = 1;
  ram[17601]  = 1;
  ram[17602]  = 1;
  ram[17603]  = 1;
  ram[17604]  = 1;
  ram[17605]  = 1;
  ram[17606]  = 1;
  ram[17607]  = 1;
  ram[17608]  = 1;
  ram[17609]  = 1;
  ram[17610]  = 1;
  ram[17611]  = 1;
  ram[17612]  = 1;
  ram[17613]  = 1;
  ram[17614]  = 1;
  ram[17615]  = 1;
  ram[17616]  = 1;
  ram[17617]  = 1;
  ram[17618]  = 1;
  ram[17619]  = 1;
  ram[17620]  = 1;
  ram[17621]  = 1;
  ram[17622]  = 1;
  ram[17623]  = 1;
  ram[17624]  = 1;
  ram[17625]  = 1;
  ram[17626]  = 1;
  ram[17627]  = 1;
  ram[17628]  = 1;
  ram[17629]  = 1;
  ram[17630]  = 1;
  ram[17631]  = 1;
  ram[17632]  = 1;
  ram[17633]  = 1;
  ram[17634]  = 1;
  ram[17635]  = 1;
  ram[17636]  = 1;
  ram[17637]  = 1;
  ram[17638]  = 1;
  ram[17639]  = 1;
  ram[17640]  = 1;
  ram[17641]  = 1;
  ram[17642]  = 1;
  ram[17643]  = 1;
  ram[17644]  = 1;
  ram[17645]  = 1;
  ram[17646]  = 1;
  ram[17647]  = 1;
  ram[17648]  = 1;
  ram[17649]  = 1;
  ram[17650]  = 1;
  ram[17651]  = 1;
  ram[17652]  = 1;
  ram[17653]  = 1;
  ram[17654]  = 1;
  ram[17655]  = 1;
  ram[17656]  = 1;
  ram[17657]  = 1;
  ram[17658]  = 1;
  ram[17659]  = 1;
  ram[17660]  = 1;
  ram[17661]  = 1;
  ram[17662]  = 1;
  ram[17663]  = 1;
  ram[17664]  = 1;
  ram[17665]  = 1;
  ram[17666]  = 1;
  ram[17667]  = 1;
  ram[17668]  = 1;
  ram[17669]  = 1;
  ram[17670]  = 1;
  ram[17671]  = 1;
  ram[17672]  = 1;
  ram[17673]  = 1;
  ram[17674]  = 1;
  ram[17675]  = 1;
  ram[17676]  = 1;
  ram[17677]  = 1;
  ram[17678]  = 1;
  ram[17679]  = 1;
  ram[17680]  = 1;
  ram[17681]  = 1;
  ram[17682]  = 1;
  ram[17683]  = 1;
  ram[17684]  = 1;
  ram[17685]  = 1;
  ram[17686]  = 1;
  ram[17687]  = 1;
  ram[17688]  = 1;
  ram[17689]  = 1;
  ram[17690]  = 1;
  ram[17691]  = 1;
  ram[17692]  = 1;
  ram[17693]  = 1;
  ram[17694]  = 1;
  ram[17695]  = 1;
  ram[17696]  = 1;
  ram[17697]  = 1;
  ram[17698]  = 1;
  ram[17699]  = 1;
  ram[17700]  = 1;
  ram[17701]  = 1;
  ram[17702]  = 1;
  ram[17703]  = 1;
  ram[17704]  = 1;
  ram[17705]  = 1;
  ram[17706]  = 1;
  ram[17707]  = 1;
  ram[17708]  = 1;
  ram[17709]  = 1;
  ram[17710]  = 1;
  ram[17711]  = 1;
  ram[17712]  = 1;
  ram[17713]  = 1;
  ram[17714]  = 1;
  ram[17715]  = 1;
  ram[17716]  = 1;
  ram[17717]  = 1;
  ram[17718]  = 1;
  ram[17719]  = 1;
  ram[17720]  = 1;
  ram[17721]  = 1;
  ram[17722]  = 1;
  ram[17723]  = 1;
  ram[17724]  = 1;
  ram[17725]  = 1;
  ram[17726]  = 1;
  ram[17727]  = 1;
  ram[17728]  = 1;
  ram[17729]  = 1;
  ram[17730]  = 1;
  ram[17731]  = 1;
  ram[17732]  = 1;
  ram[17733]  = 1;
  ram[17734]  = 1;
  ram[17735]  = 1;
  ram[17736]  = 1;
  ram[17737]  = 1;
  ram[17738]  = 1;
  ram[17739]  = 1;
  ram[17740]  = 1;
  ram[17741]  = 1;
  ram[17742]  = 1;
  ram[17743]  = 1;
  ram[17744]  = 1;
  ram[17745]  = 1;
  ram[17746]  = 1;
  ram[17747]  = 1;
  ram[17748]  = 1;
  ram[17749]  = 1;
  ram[17750]  = 1;
  ram[17751]  = 1;
  ram[17752]  = 1;
  ram[17753]  = 1;
  ram[17754]  = 1;
  ram[17755]  = 1;
  ram[17756]  = 1;
  ram[17757]  = 1;
  ram[17758]  = 1;
  ram[17759]  = 1;
  ram[17760]  = 1;
  ram[17761]  = 1;
  ram[17762]  = 1;
  ram[17763]  = 1;
  ram[17764]  = 1;
  ram[17765]  = 1;
  ram[17766]  = 1;
  ram[17767]  = 1;
  ram[17768]  = 1;
  ram[17769]  = 1;
  ram[17770]  = 1;
  ram[17771]  = 1;
  ram[17772]  = 1;
  ram[17773]  = 1;
  ram[17774]  = 1;
  ram[17775]  = 1;
  ram[17776]  = 1;
  ram[17777]  = 1;
  ram[17778]  = 1;
  ram[17779]  = 1;
  ram[17780]  = 1;
  ram[17781]  = 1;
  ram[17782]  = 1;
  ram[17783]  = 1;
  ram[17784]  = 1;
  ram[17785]  = 1;
  ram[17786]  = 1;
  ram[17787]  = 1;
  ram[17788]  = 1;
  ram[17789]  = 1;
  ram[17790]  = 1;
  ram[17791]  = 1;
  ram[17792]  = 1;
  ram[17793]  = 1;
  ram[17794]  = 1;
  ram[17795]  = 1;
  ram[17796]  = 1;
  ram[17797]  = 1;
  ram[17798]  = 1;
  ram[17799]  = 1;
  ram[17800]  = 1;
  ram[17801]  = 1;
  ram[17802]  = 1;
  ram[17803]  = 1;
  ram[17804]  = 1;
  ram[17805]  = 1;
  ram[17806]  = 1;
  ram[17807]  = 1;
  ram[17808]  = 1;
  ram[17809]  = 1;
  ram[17810]  = 1;
  ram[17811]  = 1;
  ram[17812]  = 1;
  ram[17813]  = 1;
  ram[17814]  = 1;
  ram[17815]  = 1;
  ram[17816]  = 1;
  ram[17817]  = 1;
  ram[17818]  = 1;
  ram[17819]  = 1;
  ram[17820]  = 1;
  ram[17821]  = 1;
  ram[17822]  = 1;
  ram[17823]  = 1;
  ram[17824]  = 1;
  ram[17825]  = 1;
  ram[17826]  = 1;
  ram[17827]  = 1;
  ram[17828]  = 1;
  ram[17829]  = 1;
  ram[17830]  = 1;
  ram[17831]  = 1;
  ram[17832]  = 1;
  ram[17833]  = 1;
  ram[17834]  = 1;
  ram[17835]  = 1;
  ram[17836]  = 1;
  ram[17837]  = 1;
  ram[17838]  = 1;
  ram[17839]  = 1;
  ram[17840]  = 1;
  ram[17841]  = 1;
  ram[17842]  = 1;
  ram[17843]  = 1;
  ram[17844]  = 1;
  ram[17845]  = 1;
  ram[17846]  = 1;
  ram[17847]  = 1;
  ram[17848]  = 1;
  ram[17849]  = 1;
  ram[17850]  = 1;
  ram[17851]  = 1;
  ram[17852]  = 1;
  ram[17853]  = 1;
  ram[17854]  = 1;
  ram[17855]  = 1;
  ram[17856]  = 1;
  ram[17857]  = 1;
  ram[17858]  = 1;
  ram[17859]  = 1;
  ram[17860]  = 1;
  ram[17861]  = 1;
  ram[17862]  = 1;
  ram[17863]  = 1;
  ram[17864]  = 1;
  ram[17865]  = 1;
  ram[17866]  = 1;
  ram[17867]  = 1;
  ram[17868]  = 1;
  ram[17869]  = 1;
  ram[17870]  = 1;
  ram[17871]  = 1;
  ram[17872]  = 1;
  ram[17873]  = 1;
  ram[17874]  = 1;
  ram[17875]  = 1;
  ram[17876]  = 1;
  ram[17877]  = 1;
  ram[17878]  = 1;
  ram[17879]  = 1;
  ram[17880]  = 1;
  ram[17881]  = 1;
  ram[17882]  = 1;
  ram[17883]  = 1;
  ram[17884]  = 1;
  ram[17885]  = 1;
  ram[17886]  = 1;
  ram[17887]  = 1;
  ram[17888]  = 1;
  ram[17889]  = 1;
  ram[17890]  = 1;
  ram[17891]  = 1;
  ram[17892]  = 1;
  ram[17893]  = 1;
  ram[17894]  = 1;
  ram[17895]  = 1;
  ram[17896]  = 1;
  ram[17897]  = 1;
  ram[17898]  = 1;
  ram[17899]  = 1;
  ram[17900]  = 1;
  ram[17901]  = 1;
  ram[17902]  = 1;
  ram[17903]  = 1;
  ram[17904]  = 1;
  ram[17905]  = 1;
  ram[17906]  = 1;
  ram[17907]  = 1;
  ram[17908]  = 1;
  ram[17909]  = 1;
  ram[17910]  = 1;
  ram[17911]  = 1;
  ram[17912]  = 1;
  ram[17913]  = 1;
  ram[17914]  = 1;
  ram[17915]  = 1;
  ram[17916]  = 1;
  ram[17917]  = 1;
  ram[17918]  = 1;
  ram[17919]  = 1;
  ram[17920]  = 1;
  ram[17921]  = 1;
  ram[17922]  = 1;
  ram[17923]  = 1;
  ram[17924]  = 1;
  ram[17925]  = 1;
  ram[17926]  = 1;
  ram[17927]  = 1;
  ram[17928]  = 1;
  ram[17929]  = 1;
  ram[17930]  = 1;
  ram[17931]  = 1;
  ram[17932]  = 1;
  ram[17933]  = 1;
  ram[17934]  = 1;
  ram[17935]  = 1;
  ram[17936]  = 1;
  ram[17937]  = 1;
  ram[17938]  = 1;
  ram[17939]  = 1;
  ram[17940]  = 1;
  ram[17941]  = 1;
  ram[17942]  = 1;
  ram[17943]  = 1;
  ram[17944]  = 1;
  ram[17945]  = 1;
  ram[17946]  = 1;
  ram[17947]  = 1;
  ram[17948]  = 1;
  ram[17949]  = 1;
  ram[17950]  = 1;
  ram[17951]  = 1;
  ram[17952]  = 1;
  ram[17953]  = 1;
  ram[17954]  = 1;
  ram[17955]  = 1;
  ram[17956]  = 1;
  ram[17957]  = 1;
  ram[17958]  = 1;
  ram[17959]  = 1;
  ram[17960]  = 1;
  ram[17961]  = 1;
  ram[17962]  = 1;
  ram[17963]  = 1;
  ram[17964]  = 1;
  ram[17965]  = 1;
  ram[17966]  = 1;
  ram[17967]  = 1;
  ram[17968]  = 1;
  ram[17969]  = 1;
  ram[17970]  = 1;
  ram[17971]  = 1;
  ram[17972]  = 1;
  ram[17973]  = 1;
  ram[17974]  = 1;
  ram[17975]  = 1;
  ram[17976]  = 1;
  ram[17977]  = 1;
  ram[17978]  = 1;
  ram[17979]  = 1;
  ram[17980]  = 1;
  ram[17981]  = 1;
  ram[17982]  = 1;
  ram[17983]  = 1;
  ram[17984]  = 1;
  ram[17985]  = 1;
  ram[17986]  = 1;
  ram[17987]  = 1;
  ram[17988]  = 1;
  ram[17989]  = 1;
  ram[17990]  = 1;
  ram[17991]  = 1;
  ram[17992]  = 1;
  ram[17993]  = 1;
  ram[17994]  = 1;
  ram[17995]  = 1;
  ram[17996]  = 1;
  ram[17997]  = 1;
  ram[17998]  = 1;
  ram[17999]  = 1;
  ram[18000]  = 1;
  ram[18001]  = 1;
  ram[18002]  = 1;
  ram[18003]  = 1;
  ram[18004]  = 1;
  ram[18005]  = 1;
  ram[18006]  = 1;
  ram[18007]  = 1;
  ram[18008]  = 1;
  ram[18009]  = 1;
  ram[18010]  = 1;
  ram[18011]  = 1;
  ram[18012]  = 1;
  ram[18013]  = 1;
  ram[18014]  = 1;
  ram[18015]  = 1;
  ram[18016]  = 1;
  ram[18017]  = 1;
  ram[18018]  = 1;
  ram[18019]  = 1;
  ram[18020]  = 1;
  ram[18021]  = 1;
  ram[18022]  = 1;
  ram[18023]  = 1;
  ram[18024]  = 1;
  ram[18025]  = 1;
  ram[18026]  = 1;
  ram[18027]  = 1;
  ram[18028]  = 1;
  ram[18029]  = 1;
  ram[18030]  = 1;
  ram[18031]  = 1;
  ram[18032]  = 1;
  ram[18033]  = 1;
  ram[18034]  = 1;
  ram[18035]  = 1;
  ram[18036]  = 1;
  ram[18037]  = 1;
  ram[18038]  = 1;
  ram[18039]  = 1;
  ram[18040]  = 1;
  ram[18041]  = 1;
  ram[18042]  = 1;
  ram[18043]  = 1;
  ram[18044]  = 1;
  ram[18045]  = 1;
  ram[18046]  = 1;
  ram[18047]  = 1;
  ram[18048]  = 1;
  ram[18049]  = 1;
  ram[18050]  = 1;
  ram[18051]  = 1;
  ram[18052]  = 1;
  ram[18053]  = 1;
  ram[18054]  = 1;
  ram[18055]  = 1;
  ram[18056]  = 1;
  ram[18057]  = 1;
  ram[18058]  = 1;
  ram[18059]  = 1;
  ram[18060]  = 1;
  ram[18061]  = 1;
  ram[18062]  = 1;
  ram[18063]  = 1;
  ram[18064]  = 1;
  ram[18065]  = 1;
  ram[18066]  = 1;
  ram[18067]  = 1;
  ram[18068]  = 1;
  ram[18069]  = 1;
  ram[18070]  = 1;
  ram[18071]  = 1;
  ram[18072]  = 1;
  ram[18073]  = 1;
  ram[18074]  = 1;
  ram[18075]  = 1;
  ram[18076]  = 1;
  ram[18077]  = 1;
  ram[18078]  = 1;
  ram[18079]  = 1;
  ram[18080]  = 1;
  ram[18081]  = 1;
  ram[18082]  = 1;
  ram[18083]  = 1;
  ram[18084]  = 1;
  ram[18085]  = 1;
  ram[18086]  = 1;
  ram[18087]  = 1;
  ram[18088]  = 1;
  ram[18089]  = 1;
  ram[18090]  = 1;
  ram[18091]  = 1;
  ram[18092]  = 1;
  ram[18093]  = 1;
  ram[18094]  = 1;
  ram[18095]  = 1;
  ram[18096]  = 1;
  ram[18097]  = 1;
  ram[18098]  = 1;
  ram[18099]  = 1;
  ram[18100]  = 1;
  ram[18101]  = 1;
  ram[18102]  = 1;
  ram[18103]  = 1;
  ram[18104]  = 1;
  ram[18105]  = 1;
  ram[18106]  = 1;
  ram[18107]  = 1;
  ram[18108]  = 1;
  ram[18109]  = 1;
  ram[18110]  = 1;
  ram[18111]  = 1;
  ram[18112]  = 1;
  ram[18113]  = 1;
  ram[18114]  = 1;
  ram[18115]  = 1;
  ram[18116]  = 1;
  ram[18117]  = 1;
  ram[18118]  = 1;
  ram[18119]  = 1;
  ram[18120]  = 1;
  ram[18121]  = 1;
  ram[18122]  = 1;
  ram[18123]  = 1;
  ram[18124]  = 1;
  ram[18125]  = 1;
  ram[18126]  = 1;
  ram[18127]  = 1;
  ram[18128]  = 1;
  ram[18129]  = 1;
  ram[18130]  = 1;
  ram[18131]  = 1;
  ram[18132]  = 1;
  ram[18133]  = 1;
  ram[18134]  = 1;
  ram[18135]  = 1;
  ram[18136]  = 1;
  ram[18137]  = 1;
  ram[18138]  = 1;
  ram[18139]  = 1;
  ram[18140]  = 1;
  ram[18141]  = 1;
  ram[18142]  = 1;
  ram[18143]  = 1;
  ram[18144]  = 1;
  ram[18145]  = 1;
  ram[18146]  = 1;
  ram[18147]  = 1;
  ram[18148]  = 1;
  ram[18149]  = 1;
  ram[18150]  = 1;
  ram[18151]  = 1;
  ram[18152]  = 1;
  ram[18153]  = 1;
  ram[18154]  = 1;
  ram[18155]  = 1;
  ram[18156]  = 1;
  ram[18157]  = 1;
  ram[18158]  = 1;
  ram[18159]  = 1;
  ram[18160]  = 1;
  ram[18161]  = 1;
  ram[18162]  = 1;
  ram[18163]  = 1;
  ram[18164]  = 1;
  ram[18165]  = 1;
  ram[18166]  = 1;
  ram[18167]  = 1;
  ram[18168]  = 1;
  ram[18169]  = 1;
  ram[18170]  = 1;
  ram[18171]  = 1;
  ram[18172]  = 1;
  ram[18173]  = 1;
  ram[18174]  = 1;
  ram[18175]  = 1;
  ram[18176]  = 1;
  ram[18177]  = 1;
  ram[18178]  = 1;
  ram[18179]  = 1;
  ram[18180]  = 1;
  ram[18181]  = 1;
  ram[18182]  = 1;
  ram[18183]  = 1;
  ram[18184]  = 1;
  ram[18185]  = 1;
  ram[18186]  = 1;
  ram[18187]  = 1;
  ram[18188]  = 1;
  ram[18189]  = 1;
  ram[18190]  = 1;
  ram[18191]  = 1;
  ram[18192]  = 1;
  ram[18193]  = 1;
  ram[18194]  = 1;
  ram[18195]  = 1;
  ram[18196]  = 1;
  ram[18197]  = 1;
  ram[18198]  = 1;
  ram[18199]  = 1;
  ram[18200]  = 1;
  ram[18201]  = 1;
  ram[18202]  = 1;
  ram[18203]  = 1;
  ram[18204]  = 1;
  ram[18205]  = 1;
  ram[18206]  = 1;
  ram[18207]  = 1;
  ram[18208]  = 1;
  ram[18209]  = 1;
  ram[18210]  = 1;
  ram[18211]  = 1;
  ram[18212]  = 1;
  ram[18213]  = 1;
  ram[18214]  = 1;
  ram[18215]  = 1;
  ram[18216]  = 1;
  ram[18217]  = 1;
  ram[18218]  = 1;
  ram[18219]  = 1;
  ram[18220]  = 1;
  ram[18221]  = 1;
  ram[18222]  = 1;
  ram[18223]  = 1;
  ram[18224]  = 1;
  ram[18225]  = 1;
  ram[18226]  = 1;
  ram[18227]  = 1;
  ram[18228]  = 1;
  ram[18229]  = 1;
  ram[18230]  = 1;
  ram[18231]  = 1;
  ram[18232]  = 1;
  ram[18233]  = 1;
  ram[18234]  = 1;
  ram[18235]  = 1;
  ram[18236]  = 1;
  ram[18237]  = 1;
  ram[18238]  = 1;
  ram[18239]  = 1;
  ram[18240]  = 1;
  ram[18241]  = 1;
  ram[18242]  = 1;
  ram[18243]  = 1;
  ram[18244]  = 1;
  ram[18245]  = 1;
  ram[18246]  = 1;
  ram[18247]  = 1;
  ram[18248]  = 1;
  ram[18249]  = 1;
  ram[18250]  = 1;
  ram[18251]  = 1;
  ram[18252]  = 1;
  ram[18253]  = 1;
  ram[18254]  = 1;
  ram[18255]  = 1;
  ram[18256]  = 1;
  ram[18257]  = 1;
  ram[18258]  = 1;
  ram[18259]  = 1;
  ram[18260]  = 1;
  ram[18261]  = 1;
  ram[18262]  = 1;
  ram[18263]  = 1;
  ram[18264]  = 1;
  ram[18265]  = 1;
  ram[18266]  = 1;
  ram[18267]  = 1;
  ram[18268]  = 1;
  ram[18269]  = 1;
  ram[18270]  = 1;
  ram[18271]  = 1;
  ram[18272]  = 1;
  ram[18273]  = 1;
  ram[18274]  = 1;
  ram[18275]  = 1;
  ram[18276]  = 1;
  ram[18277]  = 1;
  ram[18278]  = 1;
  ram[18279]  = 1;
  ram[18280]  = 1;
  ram[18281]  = 1;
  ram[18282]  = 1;
  ram[18283]  = 1;
  ram[18284]  = 1;
  ram[18285]  = 1;
  ram[18286]  = 1;
  ram[18287]  = 1;
  ram[18288]  = 1;
  ram[18289]  = 1;
  ram[18290]  = 1;
  ram[18291]  = 1;
  ram[18292]  = 1;
  ram[18293]  = 1;
  ram[18294]  = 1;
  ram[18295]  = 1;
  ram[18296]  = 1;
  ram[18297]  = 1;
  ram[18298]  = 1;
  ram[18299]  = 1;
  ram[18300]  = 1;
  ram[18301]  = 1;
  ram[18302]  = 1;
  ram[18303]  = 1;
  ram[18304]  = 1;
  ram[18305]  = 1;
  ram[18306]  = 1;
  ram[18307]  = 1;
  ram[18308]  = 1;
  ram[18309]  = 1;
  ram[18310]  = 1;
  ram[18311]  = 1;
  ram[18312]  = 1;
  ram[18313]  = 1;
  ram[18314]  = 1;
  ram[18315]  = 1;
  ram[18316]  = 1;
  ram[18317]  = 1;
  ram[18318]  = 1;
  ram[18319]  = 1;
  ram[18320]  = 1;
  ram[18321]  = 1;
  ram[18322]  = 1;
  ram[18323]  = 1;
  ram[18324]  = 1;
  ram[18325]  = 1;
  ram[18326]  = 1;
  ram[18327]  = 1;
  ram[18328]  = 1;
  ram[18329]  = 1;
  ram[18330]  = 1;
  ram[18331]  = 1;
  ram[18332]  = 1;
  ram[18333]  = 1;
  ram[18334]  = 1;
  ram[18335]  = 1;
  ram[18336]  = 1;
  ram[18337]  = 1;
  ram[18338]  = 1;
  ram[18339]  = 1;
  ram[18340]  = 1;
  ram[18341]  = 1;
  ram[18342]  = 1;
  ram[18343]  = 1;
  ram[18344]  = 1;
  ram[18345]  = 1;
  ram[18346]  = 1;
  ram[18347]  = 1;
  ram[18348]  = 1;
  ram[18349]  = 1;
  ram[18350]  = 1;
  ram[18351]  = 1;
  ram[18352]  = 1;
  ram[18353]  = 1;
  ram[18354]  = 1;
  ram[18355]  = 1;
  ram[18356]  = 1;
  ram[18357]  = 1;
  ram[18358]  = 1;
  ram[18359]  = 1;
  ram[18360]  = 1;
  ram[18361]  = 1;
  ram[18362]  = 1;
  ram[18363]  = 1;
  ram[18364]  = 1;
  ram[18365]  = 1;
  ram[18366]  = 1;
  ram[18367]  = 1;
  ram[18368]  = 1;
  ram[18369]  = 1;
  ram[18370]  = 1;
  ram[18371]  = 1;
  ram[18372]  = 1;
  ram[18373]  = 1;
  ram[18374]  = 1;
  ram[18375]  = 1;
  ram[18376]  = 1;
  ram[18377]  = 1;
  ram[18378]  = 1;
  ram[18379]  = 1;
  ram[18380]  = 1;
  ram[18381]  = 1;
  ram[18382]  = 1;
  ram[18383]  = 1;
  ram[18384]  = 1;
  ram[18385]  = 1;
  ram[18386]  = 1;
  ram[18387]  = 1;
  ram[18388]  = 1;
  ram[18389]  = 1;
  ram[18390]  = 1;
  ram[18391]  = 1;
  ram[18392]  = 1;
  ram[18393]  = 1;
  ram[18394]  = 1;
  ram[18395]  = 1;
  ram[18396]  = 1;
  ram[18397]  = 1;
  ram[18398]  = 1;
  ram[18399]  = 1;
  ram[18400]  = 1;
  ram[18401]  = 1;
  ram[18402]  = 1;
  ram[18403]  = 1;
  ram[18404]  = 1;
  ram[18405]  = 1;
  ram[18406]  = 1;
  ram[18407]  = 1;
  ram[18408]  = 1;
  ram[18409]  = 1;
  ram[18410]  = 1;
  ram[18411]  = 1;
  ram[18412]  = 1;
  ram[18413]  = 1;
  ram[18414]  = 1;
  ram[18415]  = 1;
  ram[18416]  = 1;
  ram[18417]  = 1;
  ram[18418]  = 1;
  ram[18419]  = 1;
  ram[18420]  = 1;
  ram[18421]  = 1;
  ram[18422]  = 1;
  ram[18423]  = 1;
  ram[18424]  = 1;
  ram[18425]  = 1;
  ram[18426]  = 1;
  ram[18427]  = 1;
  ram[18428]  = 1;
  ram[18429]  = 1;
  ram[18430]  = 1;
  ram[18431]  = 1;
  ram[18432]  = 1;
  ram[18433]  = 1;
  ram[18434]  = 1;
  ram[18435]  = 1;
  ram[18436]  = 1;
  ram[18437]  = 1;
  ram[18438]  = 1;
  ram[18439]  = 1;
  ram[18440]  = 1;
  ram[18441]  = 1;
  ram[18442]  = 1;
  ram[18443]  = 1;
  ram[18444]  = 1;
  ram[18445]  = 1;
  ram[18446]  = 1;
  ram[18447]  = 1;
  ram[18448]  = 1;
  ram[18449]  = 1;
  ram[18450]  = 1;
  ram[18451]  = 1;
  ram[18452]  = 1;
  ram[18453]  = 1;
  ram[18454]  = 1;
  ram[18455]  = 1;
  ram[18456]  = 1;
  ram[18457]  = 1;
  ram[18458]  = 1;
  ram[18459]  = 1;
  ram[18460]  = 1;
  ram[18461]  = 1;
  ram[18462]  = 1;
  ram[18463]  = 1;
  ram[18464]  = 1;
  ram[18465]  = 1;
  ram[18466]  = 1;
  ram[18467]  = 1;
  ram[18468]  = 1;
  ram[18469]  = 1;
  ram[18470]  = 1;
  ram[18471]  = 1;
  ram[18472]  = 1;
  ram[18473]  = 1;
  ram[18474]  = 1;
  ram[18475]  = 1;
  ram[18476]  = 1;
  ram[18477]  = 1;
  ram[18478]  = 1;
  ram[18479]  = 1;
  ram[18480]  = 1;
  ram[18481]  = 1;
  ram[18482]  = 1;
  ram[18483]  = 1;
  ram[18484]  = 1;
  ram[18485]  = 1;
  ram[18486]  = 1;
  ram[18487]  = 1;
  ram[18488]  = 1;
  ram[18489]  = 1;
  ram[18490]  = 1;
  ram[18491]  = 1;
  ram[18492]  = 1;
  ram[18493]  = 1;
  ram[18494]  = 1;
  ram[18495]  = 1;
  ram[18496]  = 1;
  ram[18497]  = 1;
  ram[18498]  = 1;
  ram[18499]  = 1;
  ram[18500]  = 1;
  ram[18501]  = 1;
  ram[18502]  = 1;
  ram[18503]  = 1;
  ram[18504]  = 1;
  ram[18505]  = 1;
  ram[18506]  = 1;
  ram[18507]  = 1;
  ram[18508]  = 1;
  ram[18509]  = 1;
  ram[18510]  = 1;
  ram[18511]  = 1;
  ram[18512]  = 1;
  ram[18513]  = 1;
  ram[18514]  = 1;
  ram[18515]  = 1;
  ram[18516]  = 1;
  ram[18517]  = 1;
  ram[18518]  = 1;
  ram[18519]  = 1;
  ram[18520]  = 1;
  ram[18521]  = 1;
  ram[18522]  = 1;
  ram[18523]  = 1;
  ram[18524]  = 1;
  ram[18525]  = 1;
  ram[18526]  = 1;
  ram[18527]  = 1;
  ram[18528]  = 1;
  ram[18529]  = 1;
  ram[18530]  = 1;
  ram[18531]  = 1;
  ram[18532]  = 1;
  ram[18533]  = 1;
  ram[18534]  = 1;
  ram[18535]  = 1;
  ram[18536]  = 1;
  ram[18537]  = 1;
  ram[18538]  = 1;
  ram[18539]  = 1;
  ram[18540]  = 1;
  ram[18541]  = 1;
  ram[18542]  = 1;
  ram[18543]  = 1;
  ram[18544]  = 1;
  ram[18545]  = 1;
  ram[18546]  = 1;
  ram[18547]  = 1;
  ram[18548]  = 1;
  ram[18549]  = 1;
  ram[18550]  = 1;
  ram[18551]  = 1;
  ram[18552]  = 1;
  ram[18553]  = 1;
  ram[18554]  = 1;
  ram[18555]  = 1;
  ram[18556]  = 1;
  ram[18557]  = 1;
  ram[18558]  = 1;
  ram[18559]  = 1;
  ram[18560]  = 1;
  ram[18561]  = 1;
  ram[18562]  = 1;
  ram[18563]  = 1;
  ram[18564]  = 1;
  ram[18565]  = 1;
  ram[18566]  = 1;
  ram[18567]  = 1;
  ram[18568]  = 1;
  ram[18569]  = 1;
  ram[18570]  = 1;
  ram[18571]  = 1;
  ram[18572]  = 1;
  ram[18573]  = 1;
  ram[18574]  = 1;
  ram[18575]  = 1;
  ram[18576]  = 1;
  ram[18577]  = 1;
  ram[18578]  = 1;
  ram[18579]  = 1;
  ram[18580]  = 1;
  ram[18581]  = 1;
  ram[18582]  = 1;
  ram[18583]  = 1;
  ram[18584]  = 1;
  ram[18585]  = 1;
  ram[18586]  = 1;
  ram[18587]  = 1;
  ram[18588]  = 1;
  ram[18589]  = 1;
  ram[18590]  = 1;
  ram[18591]  = 1;
  ram[18592]  = 1;
  ram[18593]  = 1;
  ram[18594]  = 1;
  ram[18595]  = 1;
  ram[18596]  = 1;
  ram[18597]  = 1;
  ram[18598]  = 1;
  ram[18599]  = 1;
  ram[18600]  = 1;
  ram[18601]  = 1;
  ram[18602]  = 1;
  ram[18603]  = 1;
  ram[18604]  = 1;
  ram[18605]  = 1;
  ram[18606]  = 1;
  ram[18607]  = 1;
  ram[18608]  = 1;
  ram[18609]  = 1;
  ram[18610]  = 1;
  ram[18611]  = 1;
  ram[18612]  = 1;
  ram[18613]  = 1;
  ram[18614]  = 1;
  ram[18615]  = 1;
  ram[18616]  = 1;
  ram[18617]  = 1;
  ram[18618]  = 1;
  ram[18619]  = 1;
  ram[18620]  = 1;
  ram[18621]  = 1;
  ram[18622]  = 1;
  ram[18623]  = 1;
  ram[18624]  = 1;
  ram[18625]  = 1;
  ram[18626]  = 1;
  ram[18627]  = 1;
  ram[18628]  = 1;
  ram[18629]  = 1;
  ram[18630]  = 1;
  ram[18631]  = 1;
  ram[18632]  = 1;
  ram[18633]  = 1;
  ram[18634]  = 1;
  ram[18635]  = 1;
  ram[18636]  = 1;
  ram[18637]  = 1;
  ram[18638]  = 1;
  ram[18639]  = 1;
  ram[18640]  = 1;
  ram[18641]  = 1;
  ram[18642]  = 1;
  ram[18643]  = 1;
  ram[18644]  = 1;
  ram[18645]  = 1;
  ram[18646]  = 1;
  ram[18647]  = 1;
  ram[18648]  = 1;
  ram[18649]  = 1;
  ram[18650]  = 1;
  ram[18651]  = 1;
  ram[18652]  = 1;
  ram[18653]  = 1;
  ram[18654]  = 1;
  ram[18655]  = 1;
  ram[18656]  = 1;
  ram[18657]  = 1;
  ram[18658]  = 1;
  ram[18659]  = 1;
  ram[18660]  = 1;
  ram[18661]  = 1;
  ram[18662]  = 1;
  ram[18663]  = 1;
  ram[18664]  = 1;
  ram[18665]  = 1;
  ram[18666]  = 1;
  ram[18667]  = 1;
  ram[18668]  = 1;
  ram[18669]  = 1;
  ram[18670]  = 1;
  ram[18671]  = 1;
  ram[18672]  = 1;
  ram[18673]  = 1;
  ram[18674]  = 1;
  ram[18675]  = 1;
  ram[18676]  = 1;
  ram[18677]  = 1;
  ram[18678]  = 1;
  ram[18679]  = 1;
  ram[18680]  = 1;
  ram[18681]  = 1;
  ram[18682]  = 1;
  ram[18683]  = 1;
  ram[18684]  = 1;
  ram[18685]  = 1;
  ram[18686]  = 1;
  ram[18687]  = 1;
  ram[18688]  = 1;
  ram[18689]  = 1;
  ram[18690]  = 1;
  ram[18691]  = 1;
  ram[18692]  = 1;
  ram[18693]  = 1;
  ram[18694]  = 1;
  ram[18695]  = 1;
  ram[18696]  = 1;
  ram[18697]  = 1;
  ram[18698]  = 1;
  ram[18699]  = 1;
  ram[18700]  = 1;
  ram[18701]  = 1;
  ram[18702]  = 1;
  ram[18703]  = 1;
  ram[18704]  = 1;
  ram[18705]  = 1;
  ram[18706]  = 1;
  ram[18707]  = 1;
  ram[18708]  = 1;
  ram[18709]  = 1;
  ram[18710]  = 1;
  ram[18711]  = 1;
  ram[18712]  = 1;
  ram[18713]  = 1;
  ram[18714]  = 1;
  ram[18715]  = 1;
  ram[18716]  = 1;
  ram[18717]  = 1;
  ram[18718]  = 1;
  ram[18719]  = 1;
  ram[18720]  = 1;
  ram[18721]  = 1;
  ram[18722]  = 1;
  ram[18723]  = 1;
  ram[18724]  = 1;
  ram[18725]  = 1;
  ram[18726]  = 1;
  ram[18727]  = 1;
  ram[18728]  = 1;
  ram[18729]  = 1;
  ram[18730]  = 1;
  ram[18731]  = 1;
  ram[18732]  = 1;
  ram[18733]  = 1;
  ram[18734]  = 1;
  ram[18735]  = 1;
  ram[18736]  = 1;
  ram[18737]  = 1;
  ram[18738]  = 1;
  ram[18739]  = 1;
  ram[18740]  = 1;
  ram[18741]  = 1;
  ram[18742]  = 1;
  ram[18743]  = 1;
  ram[18744]  = 1;
  ram[18745]  = 1;
  ram[18746]  = 1;
  ram[18747]  = 1;
  ram[18748]  = 1;
  ram[18749]  = 1;
  ram[18750]  = 1;
  ram[18751]  = 1;
  ram[18752]  = 1;
  ram[18753]  = 1;
  ram[18754]  = 1;
  ram[18755]  = 1;
  ram[18756]  = 1;
  ram[18757]  = 1;
  ram[18758]  = 1;
  ram[18759]  = 1;
  ram[18760]  = 1;
  ram[18761]  = 1;
  ram[18762]  = 1;
  ram[18763]  = 1;
  ram[18764]  = 1;
  ram[18765]  = 1;
  ram[18766]  = 1;
  ram[18767]  = 1;
  ram[18768]  = 1;
  ram[18769]  = 1;
  ram[18770]  = 1;
  ram[18771]  = 1;
  ram[18772]  = 1;
  ram[18773]  = 1;
  ram[18774]  = 1;
  ram[18775]  = 1;
  ram[18776]  = 1;
  ram[18777]  = 1;
  ram[18778]  = 1;
  ram[18779]  = 1;
  ram[18780]  = 1;
  ram[18781]  = 1;
  ram[18782]  = 1;
  ram[18783]  = 1;
  ram[18784]  = 1;
  ram[18785]  = 1;
  ram[18786]  = 1;
  ram[18787]  = 1;
  ram[18788]  = 1;
  ram[18789]  = 1;
  ram[18790]  = 1;
  ram[18791]  = 1;
  ram[18792]  = 1;
  ram[18793]  = 1;
  ram[18794]  = 1;
  ram[18795]  = 1;
  ram[18796]  = 1;
  ram[18797]  = 1;
  ram[18798]  = 1;
  ram[18799]  = 1;
  ram[18800]  = 1;
  ram[18801]  = 1;
  ram[18802]  = 1;
  ram[18803]  = 1;
  ram[18804]  = 1;
  ram[18805]  = 1;
  ram[18806]  = 1;
  ram[18807]  = 1;
  ram[18808]  = 1;
  ram[18809]  = 1;
  ram[18810]  = 1;
  ram[18811]  = 1;
  ram[18812]  = 1;
  ram[18813]  = 1;
  ram[18814]  = 1;
  ram[18815]  = 1;
  ram[18816]  = 1;
  ram[18817]  = 1;
  ram[18818]  = 1;
  ram[18819]  = 1;
  ram[18820]  = 1;
  ram[18821]  = 1;
  ram[18822]  = 1;
  ram[18823]  = 1;
  ram[18824]  = 1;
  ram[18825]  = 1;
  ram[18826]  = 1;
  ram[18827]  = 1;
  ram[18828]  = 1;
  ram[18829]  = 1;
  ram[18830]  = 1;
  ram[18831]  = 1;
  ram[18832]  = 1;
  ram[18833]  = 1;
  ram[18834]  = 1;
  ram[18835]  = 1;
  ram[18836]  = 1;
  ram[18837]  = 1;
  ram[18838]  = 1;
  ram[18839]  = 1;
  ram[18840]  = 1;
  ram[18841]  = 1;
  ram[18842]  = 1;
  ram[18843]  = 1;
  ram[18844]  = 1;
  ram[18845]  = 1;
  ram[18846]  = 1;
  ram[18847]  = 1;
  ram[18848]  = 1;
  ram[18849]  = 1;
  ram[18850]  = 1;
  ram[18851]  = 1;
  ram[18852]  = 1;
  ram[18853]  = 1;
  ram[18854]  = 1;
  ram[18855]  = 1;
  ram[18856]  = 1;
  ram[18857]  = 1;
  ram[18858]  = 1;
  ram[18859]  = 1;
  ram[18860]  = 1;
  ram[18861]  = 1;
  ram[18862]  = 1;
  ram[18863]  = 1;
  ram[18864]  = 1;
  ram[18865]  = 1;
  ram[18866]  = 1;
  ram[18867]  = 1;
  ram[18868]  = 1;
  ram[18869]  = 1;
  ram[18870]  = 1;
  ram[18871]  = 1;
  ram[18872]  = 1;
  ram[18873]  = 1;
  ram[18874]  = 1;
  ram[18875]  = 1;
  ram[18876]  = 1;
  ram[18877]  = 1;
  ram[18878]  = 1;
  ram[18879]  = 1;
  ram[18880]  = 1;
  ram[18881]  = 1;
  ram[18882]  = 1;
  ram[18883]  = 1;
  ram[18884]  = 1;
  ram[18885]  = 1;
  ram[18886]  = 1;
  ram[18887]  = 1;
  ram[18888]  = 1;
  ram[18889]  = 1;
  ram[18890]  = 1;
  ram[18891]  = 1;
  ram[18892]  = 1;
  ram[18893]  = 1;
  ram[18894]  = 1;
  ram[18895]  = 1;
  ram[18896]  = 1;
  ram[18897]  = 1;
  ram[18898]  = 1;
  ram[18899]  = 1;
  ram[18900]  = 1;
  ram[18901]  = 1;
  ram[18902]  = 1;
  ram[18903]  = 1;
  ram[18904]  = 1;
  ram[18905]  = 1;
  ram[18906]  = 1;
  ram[18907]  = 1;
  ram[18908]  = 1;
  ram[18909]  = 1;
  ram[18910]  = 1;
  ram[18911]  = 1;
  ram[18912]  = 1;
  ram[18913]  = 1;
  ram[18914]  = 1;
  ram[18915]  = 1;
  ram[18916]  = 1;
  ram[18917]  = 1;
  ram[18918]  = 1;
  ram[18919]  = 1;
  ram[18920]  = 1;
  ram[18921]  = 1;
  ram[18922]  = 1;
  ram[18923]  = 1;
  ram[18924]  = 1;
  ram[18925]  = 1;
  ram[18926]  = 1;
  ram[18927]  = 1;
  ram[18928]  = 1;
  ram[18929]  = 1;
  ram[18930]  = 1;
  ram[18931]  = 1;
  ram[18932]  = 1;
  ram[18933]  = 1;
  ram[18934]  = 1;
  ram[18935]  = 1;
  ram[18936]  = 1;
  ram[18937]  = 1;
  ram[18938]  = 1;
  ram[18939]  = 1;
  ram[18940]  = 1;
  ram[18941]  = 1;
  ram[18942]  = 1;
  ram[18943]  = 1;
  ram[18944]  = 1;
  ram[18945]  = 1;
  ram[18946]  = 1;
  ram[18947]  = 1;
  ram[18948]  = 1;
  ram[18949]  = 1;
  ram[18950]  = 1;
  ram[18951]  = 1;
  ram[18952]  = 1;
  ram[18953]  = 1;
  ram[18954]  = 1;
  ram[18955]  = 1;
  ram[18956]  = 1;
  ram[18957]  = 1;
  ram[18958]  = 1;
  ram[18959]  = 1;
  ram[18960]  = 1;
  ram[18961]  = 1;
  ram[18962]  = 1;
  ram[18963]  = 1;
  ram[18964]  = 1;
  ram[18965]  = 1;
  ram[18966]  = 1;
  ram[18967]  = 1;
  ram[18968]  = 1;
  ram[18969]  = 1;
  ram[18970]  = 1;
  ram[18971]  = 1;
  ram[18972]  = 1;
  ram[18973]  = 1;
  ram[18974]  = 1;
  ram[18975]  = 1;
  ram[18976]  = 1;
  ram[18977]  = 1;
  ram[18978]  = 1;
  ram[18979]  = 1;
  ram[18980]  = 1;
  ram[18981]  = 1;
  ram[18982]  = 1;
  ram[18983]  = 1;
  ram[18984]  = 1;
  ram[18985]  = 1;
  ram[18986]  = 1;
  ram[18987]  = 1;
  ram[18988]  = 1;
  ram[18989]  = 1;
  ram[18990]  = 1;
  ram[18991]  = 1;
  ram[18992]  = 1;
  ram[18993]  = 1;
  ram[18994]  = 1;
  ram[18995]  = 1;
  ram[18996]  = 1;
  ram[18997]  = 1;
  ram[18998]  = 1;
  ram[18999]  = 1;
  ram[19000]  = 1;
  ram[19001]  = 1;
  ram[19002]  = 1;
  ram[19003]  = 1;
  ram[19004]  = 1;
  ram[19005]  = 1;
  ram[19006]  = 1;
  ram[19007]  = 1;
  ram[19008]  = 1;
  ram[19009]  = 1;
  ram[19010]  = 1;
  ram[19011]  = 1;
  ram[19012]  = 1;
  ram[19013]  = 1;
  ram[19014]  = 1;
  ram[19015]  = 1;
  ram[19016]  = 1;
  ram[19017]  = 1;
  ram[19018]  = 1;
  ram[19019]  = 1;
  ram[19020]  = 1;
  ram[19021]  = 1;
  ram[19022]  = 1;
  ram[19023]  = 1;
  ram[19024]  = 1;
  ram[19025]  = 1;
  ram[19026]  = 1;
  ram[19027]  = 1;
  ram[19028]  = 1;
  ram[19029]  = 1;
  ram[19030]  = 1;
  ram[19031]  = 1;
  ram[19032]  = 1;
  ram[19033]  = 1;
  ram[19034]  = 1;
  ram[19035]  = 1;
  ram[19036]  = 1;
  ram[19037]  = 1;
  ram[19038]  = 1;
  ram[19039]  = 1;
  ram[19040]  = 1;
  ram[19041]  = 1;
  ram[19042]  = 1;
  ram[19043]  = 1;
  ram[19044]  = 1;
  ram[19045]  = 1;
  ram[19046]  = 1;
  ram[19047]  = 1;
  ram[19048]  = 1;
  ram[19049]  = 1;
  ram[19050]  = 1;
  ram[19051]  = 1;
  ram[19052]  = 1;
  ram[19053]  = 1;
  ram[19054]  = 1;
  ram[19055]  = 1;
  ram[19056]  = 1;
  ram[19057]  = 1;
  ram[19058]  = 1;
  ram[19059]  = 1;
  ram[19060]  = 1;
  ram[19061]  = 1;
  ram[19062]  = 1;
  ram[19063]  = 1;
  ram[19064]  = 1;
  ram[19065]  = 1;
  ram[19066]  = 1;
  ram[19067]  = 1;
  ram[19068]  = 1;
  ram[19069]  = 1;
  ram[19070]  = 1;
  ram[19071]  = 1;
  ram[19072]  = 1;
  ram[19073]  = 1;
  ram[19074]  = 1;
  ram[19075]  = 1;
  ram[19076]  = 1;
  ram[19077]  = 1;
  ram[19078]  = 1;
  ram[19079]  = 1;
  ram[19080]  = 1;
  ram[19081]  = 1;
  ram[19082]  = 1;
  ram[19083]  = 1;
  ram[19084]  = 1;
  ram[19085]  = 1;
  ram[19086]  = 1;
  ram[19087]  = 1;
  ram[19088]  = 1;
  ram[19089]  = 1;
  ram[19090]  = 1;
  ram[19091]  = 1;
  ram[19092]  = 1;
  ram[19093]  = 1;
  ram[19094]  = 1;
  ram[19095]  = 1;
  ram[19096]  = 1;
  ram[19097]  = 1;
  ram[19098]  = 1;
  ram[19099]  = 1;
  ram[19100]  = 1;
  ram[19101]  = 1;
  ram[19102]  = 1;
  ram[19103]  = 1;
  ram[19104]  = 1;
  ram[19105]  = 1;
  ram[19106]  = 1;
  ram[19107]  = 1;
  ram[19108]  = 1;
  ram[19109]  = 1;
  ram[19110]  = 1;
  ram[19111]  = 1;
  ram[19112]  = 1;
  ram[19113]  = 1;
  ram[19114]  = 1;
  ram[19115]  = 1;
  ram[19116]  = 1;
  ram[19117]  = 1;
  ram[19118]  = 1;
  ram[19119]  = 1;
  ram[19120]  = 1;
  ram[19121]  = 1;
  ram[19122]  = 1;
  ram[19123]  = 1;
  ram[19124]  = 1;
  ram[19125]  = 1;
  ram[19126]  = 1;
  ram[19127]  = 1;
  ram[19128]  = 1;
  ram[19129]  = 1;
  ram[19130]  = 1;
  ram[19131]  = 1;
  ram[19132]  = 1;
  ram[19133]  = 1;
  ram[19134]  = 1;
  ram[19135]  = 1;
  ram[19136]  = 1;
  ram[19137]  = 1;
  ram[19138]  = 1;
  ram[19139]  = 1;
  ram[19140]  = 1;
  ram[19141]  = 1;
  ram[19142]  = 1;
  ram[19143]  = 1;
  ram[19144]  = 1;
  ram[19145]  = 1;
  ram[19146]  = 1;
  ram[19147]  = 1;
  ram[19148]  = 1;
  ram[19149]  = 1;
  ram[19150]  = 1;
  ram[19151]  = 1;
  ram[19152]  = 1;
  ram[19153]  = 1;
  ram[19154]  = 1;
  ram[19155]  = 1;
  ram[19156]  = 1;
  ram[19157]  = 1;
  ram[19158]  = 1;
  ram[19159]  = 1;
  ram[19160]  = 1;
  ram[19161]  = 1;
  ram[19162]  = 1;
  ram[19163]  = 1;
  ram[19164]  = 1;
  ram[19165]  = 1;
  ram[19166]  = 1;
  ram[19167]  = 1;
  ram[19168]  = 1;
  ram[19169]  = 1;
  ram[19170]  = 1;
  ram[19171]  = 1;
  ram[19172]  = 1;
  ram[19173]  = 1;
  ram[19174]  = 1;
  ram[19175]  = 1;
  ram[19176]  = 1;
  ram[19177]  = 1;
  ram[19178]  = 1;
  ram[19179]  = 1;
  ram[19180]  = 1;
  ram[19181]  = 1;
  ram[19182]  = 1;
  ram[19183]  = 1;
  ram[19184]  = 1;
  ram[19185]  = 1;
  ram[19186]  = 1;
  ram[19187]  = 1;
  ram[19188]  = 1;
  ram[19189]  = 1;
  ram[19190]  = 1;
  ram[19191]  = 1;
  ram[19192]  = 1;
  ram[19193]  = 1;
  ram[19194]  = 1;
  ram[19195]  = 1;
  ram[19196]  = 1;
  ram[19197]  = 1;
  ram[19198]  = 1;
  ram[19199]  = 1;
  ram[19200]  = 1;
  ram[19201]  = 1;
  ram[19202]  = 1;
  ram[19203]  = 1;
  ram[19204]  = 1;
  ram[19205]  = 1;
  ram[19206]  = 1;
  ram[19207]  = 1;
  ram[19208]  = 1;
  ram[19209]  = 1;
  ram[19210]  = 1;
  ram[19211]  = 1;
  ram[19212]  = 1;
  ram[19213]  = 1;
  ram[19214]  = 1;
  ram[19215]  = 1;
  ram[19216]  = 1;
  ram[19217]  = 1;
  ram[19218]  = 1;
  ram[19219]  = 1;
  ram[19220]  = 1;
  ram[19221]  = 1;
  ram[19222]  = 1;
  ram[19223]  = 1;
  ram[19224]  = 1;
  ram[19225]  = 1;
  ram[19226]  = 1;
  ram[19227]  = 1;
  ram[19228]  = 1;
  ram[19229]  = 1;
  ram[19230]  = 1;
  ram[19231]  = 1;
  ram[19232]  = 1;
  ram[19233]  = 1;
  ram[19234]  = 1;
  ram[19235]  = 1;
  ram[19236]  = 1;
  ram[19237]  = 1;
  ram[19238]  = 1;
  ram[19239]  = 1;
  ram[19240]  = 1;
  ram[19241]  = 1;
  ram[19242]  = 1;
  ram[19243]  = 1;
  ram[19244]  = 1;
  ram[19245]  = 1;
  ram[19246]  = 1;
  ram[19247]  = 1;
  ram[19248]  = 1;
  ram[19249]  = 1;
  ram[19250]  = 1;
  ram[19251]  = 1;
  ram[19252]  = 1;
  ram[19253]  = 1;
  ram[19254]  = 1;
  ram[19255]  = 1;
  ram[19256]  = 1;
  ram[19257]  = 1;
  ram[19258]  = 1;
  ram[19259]  = 1;
  ram[19260]  = 1;
  ram[19261]  = 1;
  ram[19262]  = 1;
  ram[19263]  = 1;
  ram[19264]  = 1;
  ram[19265]  = 1;
  ram[19266]  = 1;
  ram[19267]  = 1;
  ram[19268]  = 1;
  ram[19269]  = 1;
  ram[19270]  = 1;
  ram[19271]  = 1;
  ram[19272]  = 1;
  ram[19273]  = 1;
  ram[19274]  = 1;
  ram[19275]  = 1;
  ram[19276]  = 1;
  ram[19277]  = 1;
  ram[19278]  = 1;
  ram[19279]  = 1;
  ram[19280]  = 1;
  ram[19281]  = 1;
  ram[19282]  = 1;
  ram[19283]  = 1;
  ram[19284]  = 1;
  ram[19285]  = 1;
  ram[19286]  = 1;
  ram[19287]  = 1;
  ram[19288]  = 1;
  ram[19289]  = 1;
  ram[19290]  = 1;
  ram[19291]  = 1;
  ram[19292]  = 1;
  ram[19293]  = 1;
  ram[19294]  = 1;
  ram[19295]  = 1;
  ram[19296]  = 1;
  ram[19297]  = 1;
  ram[19298]  = 1;
  ram[19299]  = 1;
  ram[19300]  = 1;
  ram[19301]  = 1;
  ram[19302]  = 1;
  ram[19303]  = 1;
  ram[19304]  = 1;
  ram[19305]  = 1;
  ram[19306]  = 1;
  ram[19307]  = 1;
  ram[19308]  = 1;
  ram[19309]  = 1;
  ram[19310]  = 1;
  ram[19311]  = 1;
  ram[19312]  = 1;
  ram[19313]  = 1;
  ram[19314]  = 1;
  ram[19315]  = 1;
  ram[19316]  = 1;
  ram[19317]  = 1;
  ram[19318]  = 1;
  ram[19319]  = 1;
  ram[19320]  = 1;
  ram[19321]  = 1;
  ram[19322]  = 1;
  ram[19323]  = 1;
  ram[19324]  = 1;
  ram[19325]  = 1;
  ram[19326]  = 1;
  ram[19327]  = 1;
  ram[19328]  = 1;
  ram[19329]  = 1;
  ram[19330]  = 1;
  ram[19331]  = 1;
  ram[19332]  = 1;
  ram[19333]  = 1;
  ram[19334]  = 1;
  ram[19335]  = 1;
  ram[19336]  = 1;
  ram[19337]  = 1;
  ram[19338]  = 1;
  ram[19339]  = 1;
  ram[19340]  = 1;
  ram[19341]  = 1;
  ram[19342]  = 1;
  ram[19343]  = 1;
  ram[19344]  = 1;
  ram[19345]  = 1;
  ram[19346]  = 1;
  ram[19347]  = 1;
  ram[19348]  = 1;
  ram[19349]  = 1;
  ram[19350]  = 1;
  ram[19351]  = 1;
  ram[19352]  = 1;
  ram[19353]  = 1;
  ram[19354]  = 1;
  ram[19355]  = 1;
  ram[19356]  = 1;
  ram[19357]  = 1;
  ram[19358]  = 1;
  ram[19359]  = 1;
  ram[19360]  = 1;
  ram[19361]  = 1;
  ram[19362]  = 1;
  ram[19363]  = 1;
  ram[19364]  = 1;
  ram[19365]  = 1;
  ram[19366]  = 1;
  ram[19367]  = 1;
  ram[19368]  = 1;
  ram[19369]  = 1;
  ram[19370]  = 1;
  ram[19371]  = 1;
  ram[19372]  = 1;
  ram[19373]  = 1;
  ram[19374]  = 1;
  ram[19375]  = 1;
  ram[19376]  = 1;
  ram[19377]  = 1;
  ram[19378]  = 1;
  ram[19379]  = 1;
  ram[19380]  = 1;
  ram[19381]  = 1;
  ram[19382]  = 1;
  ram[19383]  = 1;
  ram[19384]  = 1;
  ram[19385]  = 1;
  ram[19386]  = 1;
  ram[19387]  = 1;
  ram[19388]  = 1;
  ram[19389]  = 1;
  ram[19390]  = 1;
  ram[19391]  = 1;
  ram[19392]  = 1;
  ram[19393]  = 1;
  ram[19394]  = 1;
  ram[19395]  = 1;
  ram[19396]  = 1;
  ram[19397]  = 1;
  ram[19398]  = 1;
  ram[19399]  = 1;
  ram[19400]  = 1;
  ram[19401]  = 1;
  ram[19402]  = 1;
  ram[19403]  = 1;
  ram[19404]  = 1;
  ram[19405]  = 1;
  ram[19406]  = 1;
  ram[19407]  = 1;
  ram[19408]  = 1;
  ram[19409]  = 1;
  ram[19410]  = 1;
  ram[19411]  = 1;
  ram[19412]  = 1;
  ram[19413]  = 1;
  ram[19414]  = 1;
  ram[19415]  = 1;
  ram[19416]  = 1;
  ram[19417]  = 1;
  ram[19418]  = 1;
  ram[19419]  = 1;
  ram[19420]  = 1;
  ram[19421]  = 1;
  ram[19422]  = 1;
  ram[19423]  = 1;
  ram[19424]  = 1;
  ram[19425]  = 1;
  ram[19426]  = 1;
  ram[19427]  = 1;
  ram[19428]  = 1;
  ram[19429]  = 1;
  ram[19430]  = 1;
  ram[19431]  = 1;
  ram[19432]  = 1;
  ram[19433]  = 1;
  ram[19434]  = 1;
  ram[19435]  = 1;
  ram[19436]  = 1;
  ram[19437]  = 1;
  ram[19438]  = 1;
  ram[19439]  = 1;
  ram[19440]  = 1;
  ram[19441]  = 1;
  ram[19442]  = 1;
  ram[19443]  = 1;
  ram[19444]  = 1;
  ram[19445]  = 1;
  ram[19446]  = 1;
  ram[19447]  = 1;
  ram[19448]  = 1;
  ram[19449]  = 1;
  ram[19450]  = 1;
  ram[19451]  = 1;
  ram[19452]  = 1;
  ram[19453]  = 1;
  ram[19454]  = 1;
  ram[19455]  = 1;
  ram[19456]  = 1;
  ram[19457]  = 1;
  ram[19458]  = 1;
  ram[19459]  = 1;
  ram[19460]  = 1;
  ram[19461]  = 1;
  ram[19462]  = 1;
  ram[19463]  = 1;
  ram[19464]  = 1;
  ram[19465]  = 1;
  ram[19466]  = 1;
  ram[19467]  = 1;
  ram[19468]  = 1;
  ram[19469]  = 1;
  ram[19470]  = 1;
  ram[19471]  = 1;
  ram[19472]  = 1;
  ram[19473]  = 1;
  ram[19474]  = 1;
  ram[19475]  = 1;
  ram[19476]  = 1;
  ram[19477]  = 1;
  ram[19478]  = 1;
  ram[19479]  = 1;
  ram[19480]  = 1;
  ram[19481]  = 1;
  ram[19482]  = 1;
  ram[19483]  = 1;
  ram[19484]  = 1;
  ram[19485]  = 1;
  ram[19486]  = 1;
  ram[19487]  = 1;
  ram[19488]  = 1;
  ram[19489]  = 1;
  ram[19490]  = 1;
  ram[19491]  = 1;
  ram[19492]  = 1;
  ram[19493]  = 1;
  ram[19494]  = 1;
  ram[19495]  = 1;
  ram[19496]  = 1;
  ram[19497]  = 1;
  ram[19498]  = 1;
  ram[19499]  = 1;
  ram[19500]  = 1;
  ram[19501]  = 1;
  ram[19502]  = 1;
  ram[19503]  = 1;
  ram[19504]  = 1;
  ram[19505]  = 1;
  ram[19506]  = 1;
  ram[19507]  = 1;
  ram[19508]  = 1;
  ram[19509]  = 1;
  ram[19510]  = 1;
  ram[19511]  = 1;
  ram[19512]  = 1;
  ram[19513]  = 1;
  ram[19514]  = 1;
  ram[19515]  = 1;
  ram[19516]  = 1;
  ram[19517]  = 1;
  ram[19518]  = 1;
  ram[19519]  = 1;
  ram[19520]  = 1;
  ram[19521]  = 1;
  ram[19522]  = 1;
  ram[19523]  = 1;
  ram[19524]  = 1;
  ram[19525]  = 1;
  ram[19526]  = 1;
  ram[19527]  = 1;
  ram[19528]  = 1;
  ram[19529]  = 1;
  ram[19530]  = 1;
  ram[19531]  = 1;
  ram[19532]  = 1;
  ram[19533]  = 1;
  ram[19534]  = 1;
  ram[19535]  = 1;
  ram[19536]  = 1;
  ram[19537]  = 1;
  ram[19538]  = 1;
  ram[19539]  = 1;
  ram[19540]  = 1;
  ram[19541]  = 1;
  ram[19542]  = 1;
  ram[19543]  = 1;
  ram[19544]  = 1;
  ram[19545]  = 1;
  ram[19546]  = 1;
  ram[19547]  = 1;
  ram[19548]  = 1;
  ram[19549]  = 1;
  ram[19550]  = 1;
  ram[19551]  = 1;
  ram[19552]  = 1;
  ram[19553]  = 1;
  ram[19554]  = 1;
  ram[19555]  = 1;
  ram[19556]  = 1;
  ram[19557]  = 1;
  ram[19558]  = 1;
  ram[19559]  = 1;
  ram[19560]  = 1;
  ram[19561]  = 1;
  ram[19562]  = 1;
  ram[19563]  = 1;
  ram[19564]  = 1;
  ram[19565]  = 1;
  ram[19566]  = 1;
  ram[19567]  = 1;
  ram[19568]  = 1;
  ram[19569]  = 1;
  ram[19570]  = 1;
  ram[19571]  = 1;
  ram[19572]  = 1;
  ram[19573]  = 1;
  ram[19574]  = 1;
  ram[19575]  = 1;
  ram[19576]  = 1;
  ram[19577]  = 1;
  ram[19578]  = 1;
  ram[19579]  = 1;
  ram[19580]  = 1;
  ram[19581]  = 1;
  ram[19582]  = 1;
  ram[19583]  = 1;
  ram[19584]  = 1;
  ram[19585]  = 1;
  ram[19586]  = 1;
  ram[19587]  = 1;
  ram[19588]  = 1;
  ram[19589]  = 1;
  ram[19590]  = 1;
  ram[19591]  = 1;
  ram[19592]  = 1;
  ram[19593]  = 1;
  ram[19594]  = 1;
  ram[19595]  = 1;
  ram[19596]  = 1;
  ram[19597]  = 1;
  ram[19598]  = 1;
  ram[19599]  = 1;
  ram[19600]  = 1;
  ram[19601]  = 1;
  ram[19602]  = 1;
  ram[19603]  = 1;
  ram[19604]  = 1;
  ram[19605]  = 1;
  ram[19606]  = 1;
  ram[19607]  = 1;
  ram[19608]  = 1;
  ram[19609]  = 1;
  ram[19610]  = 1;
  ram[19611]  = 1;
  ram[19612]  = 1;
  ram[19613]  = 1;
  ram[19614]  = 1;
  ram[19615]  = 1;
  ram[19616]  = 1;
  ram[19617]  = 1;
  ram[19618]  = 1;
  ram[19619]  = 1;
  ram[19620]  = 1;
  ram[19621]  = 1;
  ram[19622]  = 1;
  ram[19623]  = 1;
  ram[19624]  = 1;
  ram[19625]  = 1;
  ram[19626]  = 1;
  ram[19627]  = 1;
  ram[19628]  = 1;
  ram[19629]  = 1;
  ram[19630]  = 1;
  ram[19631]  = 1;
  ram[19632]  = 1;
  ram[19633]  = 1;
  ram[19634]  = 1;
  ram[19635]  = 1;
  ram[19636]  = 1;
  ram[19637]  = 1;
  ram[19638]  = 1;
  ram[19639]  = 1;
  ram[19640]  = 1;
  ram[19641]  = 1;
  ram[19642]  = 1;
  ram[19643]  = 1;
  ram[19644]  = 1;
  ram[19645]  = 1;
  ram[19646]  = 1;
  ram[19647]  = 1;
  ram[19648]  = 1;
  ram[19649]  = 1;
  ram[19650]  = 1;
  ram[19651]  = 1;
  ram[19652]  = 1;
  ram[19653]  = 1;
  ram[19654]  = 1;
  ram[19655]  = 1;
  ram[19656]  = 1;
  ram[19657]  = 1;
  ram[19658]  = 1;
  ram[19659]  = 1;
  ram[19660]  = 1;
  ram[19661]  = 1;
  ram[19662]  = 1;
  ram[19663]  = 1;
  ram[19664]  = 1;
  ram[19665]  = 1;
  ram[19666]  = 1;
  ram[19667]  = 1;
  ram[19668]  = 1;
  ram[19669]  = 1;
  ram[19670]  = 1;
  ram[19671]  = 1;
  ram[19672]  = 1;
  ram[19673]  = 1;
  ram[19674]  = 1;
  ram[19675]  = 1;
  ram[19676]  = 1;
  ram[19677]  = 1;
  ram[19678]  = 1;
  ram[19679]  = 1;
  ram[19680]  = 1;
  ram[19681]  = 1;
  ram[19682]  = 1;
  ram[19683]  = 1;
  ram[19684]  = 1;
  ram[19685]  = 1;
  ram[19686]  = 1;
  ram[19687]  = 1;
  ram[19688]  = 1;
  ram[19689]  = 1;
  ram[19690]  = 1;
  ram[19691]  = 1;
  ram[19692]  = 1;
  ram[19693]  = 1;
  ram[19694]  = 1;
  ram[19695]  = 1;
  ram[19696]  = 1;
  ram[19697]  = 1;
  ram[19698]  = 1;
  ram[19699]  = 1;
  ram[19700]  = 1;
  ram[19701]  = 1;
  ram[19702]  = 1;
  ram[19703]  = 1;
  ram[19704]  = 1;
  ram[19705]  = 1;
  ram[19706]  = 1;
  ram[19707]  = 1;
  ram[19708]  = 1;
  ram[19709]  = 1;
  ram[19710]  = 1;
  ram[19711]  = 1;
  ram[19712]  = 1;
  ram[19713]  = 1;
  ram[19714]  = 1;
  ram[19715]  = 1;
  ram[19716]  = 1;
  ram[19717]  = 1;
  ram[19718]  = 1;
  ram[19719]  = 1;
  ram[19720]  = 1;
  ram[19721]  = 1;
  ram[19722]  = 1;
  ram[19723]  = 1;
  ram[19724]  = 1;
  ram[19725]  = 1;
  ram[19726]  = 1;
  ram[19727]  = 1;
  ram[19728]  = 1;
  ram[19729]  = 1;
  ram[19730]  = 1;
  ram[19731]  = 1;
  ram[19732]  = 1;
  ram[19733]  = 1;
  ram[19734]  = 1;
  ram[19735]  = 1;
  ram[19736]  = 1;
  ram[19737]  = 1;
  ram[19738]  = 1;
  ram[19739]  = 1;
  ram[19740]  = 1;
  ram[19741]  = 1;
  ram[19742]  = 1;
  ram[19743]  = 1;
  ram[19744]  = 1;
  ram[19745]  = 1;
  ram[19746]  = 1;
  ram[19747]  = 1;
  ram[19748]  = 1;
  ram[19749]  = 1;
  ram[19750]  = 1;
  ram[19751]  = 1;
  ram[19752]  = 1;
  ram[19753]  = 1;
  ram[19754]  = 1;
  ram[19755]  = 1;
  ram[19756]  = 1;
  ram[19757]  = 1;
  ram[19758]  = 1;
  ram[19759]  = 1;
  ram[19760]  = 1;
  ram[19761]  = 1;
  ram[19762]  = 1;
  ram[19763]  = 1;
  ram[19764]  = 1;
  ram[19765]  = 1;
  ram[19766]  = 1;
  ram[19767]  = 1;
  ram[19768]  = 1;
  ram[19769]  = 1;
  ram[19770]  = 1;
  ram[19771]  = 1;
  ram[19772]  = 1;
  ram[19773]  = 1;
  ram[19774]  = 1;
  ram[19775]  = 1;
  ram[19776]  = 1;
  ram[19777]  = 1;
  ram[19778]  = 1;
  ram[19779]  = 1;
  ram[19780]  = 1;
  ram[19781]  = 1;
  ram[19782]  = 1;
  ram[19783]  = 1;
  ram[19784]  = 1;
  ram[19785]  = 1;
  ram[19786]  = 1;
  ram[19787]  = 1;
  ram[19788]  = 1;
  ram[19789]  = 1;
  ram[19790]  = 1;
  ram[19791]  = 1;
  ram[19792]  = 1;
  ram[19793]  = 1;
  ram[19794]  = 1;
  ram[19795]  = 1;
  ram[19796]  = 1;
  ram[19797]  = 1;
  ram[19798]  = 1;
  ram[19799]  = 1;
  ram[19800]  = 1;
  ram[19801]  = 1;
  ram[19802]  = 1;
  ram[19803]  = 1;
  ram[19804]  = 1;
  ram[19805]  = 1;
  ram[19806]  = 1;
  ram[19807]  = 1;
  ram[19808]  = 1;
  ram[19809]  = 1;
  ram[19810]  = 1;
  ram[19811]  = 1;
  ram[19812]  = 1;
  ram[19813]  = 1;
  ram[19814]  = 1;
  ram[19815]  = 1;
  ram[19816]  = 1;
  ram[19817]  = 1;
  ram[19818]  = 1;
  ram[19819]  = 1;
  ram[19820]  = 1;
  ram[19821]  = 1;
  ram[19822]  = 1;
  ram[19823]  = 1;
  ram[19824]  = 1;
  ram[19825]  = 1;
  ram[19826]  = 1;
  ram[19827]  = 1;
  ram[19828]  = 1;
  ram[19829]  = 1;
  ram[19830]  = 1;
  ram[19831]  = 1;
  ram[19832]  = 1;
  ram[19833]  = 1;
  ram[19834]  = 1;
  ram[19835]  = 1;
  ram[19836]  = 1;
  ram[19837]  = 1;
  ram[19838]  = 1;
  ram[19839]  = 1;
  ram[19840]  = 1;
  ram[19841]  = 1;
  ram[19842]  = 1;
  ram[19843]  = 1;
  ram[19844]  = 1;
  ram[19845]  = 1;
  ram[19846]  = 1;
  ram[19847]  = 1;
  ram[19848]  = 1;
  ram[19849]  = 1;
  ram[19850]  = 1;
  ram[19851]  = 1;
  ram[19852]  = 1;
  ram[19853]  = 1;
  ram[19854]  = 1;
  ram[19855]  = 1;
  ram[19856]  = 1;
  ram[19857]  = 1;
  ram[19858]  = 1;
  ram[19859]  = 1;
  ram[19860]  = 1;
  ram[19861]  = 1;
  ram[19862]  = 1;
  ram[19863]  = 1;
  ram[19864]  = 1;
  ram[19865]  = 1;
  ram[19866]  = 1;
  ram[19867]  = 1;
  ram[19868]  = 1;
  ram[19869]  = 1;
  ram[19870]  = 1;
  ram[19871]  = 1;
  ram[19872]  = 1;
  ram[19873]  = 1;
  ram[19874]  = 1;
  ram[19875]  = 1;
  ram[19876]  = 1;
  ram[19877]  = 1;
  ram[19878]  = 1;
  ram[19879]  = 1;
  ram[19880]  = 1;
  ram[19881]  = 1;
  ram[19882]  = 1;
  ram[19883]  = 1;
  ram[19884]  = 1;
  ram[19885]  = 1;
  ram[19886]  = 1;
  ram[19887]  = 1;
  ram[19888]  = 1;
  ram[19889]  = 1;
  ram[19890]  = 1;
  ram[19891]  = 1;
  ram[19892]  = 1;
  ram[19893]  = 1;
  ram[19894]  = 1;
  ram[19895]  = 1;
  ram[19896]  = 1;
  ram[19897]  = 1;
  ram[19898]  = 1;
  ram[19899]  = 1;
  ram[19900]  = 1;
  ram[19901]  = 1;
  ram[19902]  = 1;
  ram[19903]  = 1;
  ram[19904]  = 1;
  ram[19905]  = 1;
  ram[19906]  = 1;
  ram[19907]  = 1;
  ram[19908]  = 1;
  ram[19909]  = 1;
  ram[19910]  = 1;
  ram[19911]  = 1;
  ram[19912]  = 1;
  ram[19913]  = 1;
  ram[19914]  = 1;
  ram[19915]  = 1;
  ram[19916]  = 1;
  ram[19917]  = 1;
  ram[19918]  = 1;
  ram[19919]  = 1;
  ram[19920]  = 1;
  ram[19921]  = 1;
  ram[19922]  = 1;
  ram[19923]  = 1;
  ram[19924]  = 1;
  ram[19925]  = 1;
  ram[19926]  = 1;
  ram[19927]  = 1;
  ram[19928]  = 1;
  ram[19929]  = 1;
  ram[19930]  = 1;
  ram[19931]  = 1;
  ram[19932]  = 1;
  ram[19933]  = 1;
  ram[19934]  = 1;
  ram[19935]  = 1;
  ram[19936]  = 1;
  ram[19937]  = 1;
  ram[19938]  = 1;
  ram[19939]  = 1;
  ram[19940]  = 1;
  ram[19941]  = 1;
  ram[19942]  = 1;
  ram[19943]  = 1;
  ram[19944]  = 1;
  ram[19945]  = 1;
  ram[19946]  = 1;
  ram[19947]  = 1;
  ram[19948]  = 1;
  ram[19949]  = 1;
  ram[19950]  = 1;
  ram[19951]  = 1;
  ram[19952]  = 1;
  ram[19953]  = 1;
  ram[19954]  = 1;
  ram[19955]  = 1;
  ram[19956]  = 1;
  ram[19957]  = 1;
  ram[19958]  = 1;
  ram[19959]  = 1;
  ram[19960]  = 1;
  ram[19961]  = 1;
  ram[19962]  = 1;
  ram[19963]  = 1;
  ram[19964]  = 1;
  ram[19965]  = 1;
  ram[19966]  = 1;
  ram[19967]  = 1;
  ram[19968]  = 1;
  ram[19969]  = 1;
  ram[19970]  = 1;
  ram[19971]  = 1;
  ram[19972]  = 1;
  ram[19973]  = 1;
  ram[19974]  = 1;
  ram[19975]  = 1;
  ram[19976]  = 1;
  ram[19977]  = 1;
  ram[19978]  = 1;
  ram[19979]  = 1;
  ram[19980]  = 1;
  ram[19981]  = 1;
  ram[19982]  = 1;
  ram[19983]  = 1;
  ram[19984]  = 1;
  ram[19985]  = 1;
  ram[19986]  = 1;
  ram[19987]  = 1;
  ram[19988]  = 1;
  ram[19989]  = 1;
  ram[19990]  = 1;
  ram[19991]  = 1;
  ram[19992]  = 1;
  ram[19993]  = 1;
  ram[19994]  = 1;
  ram[19995]  = 1;
  ram[19996]  = 1;
  ram[19997]  = 1;
  ram[19998]  = 1;
  ram[19999]  = 1;
end

always @(posedge clock) begin
  dout <= ram[address];
end

endmodule
